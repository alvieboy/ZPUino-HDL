library IEEE;
use IEEE.std_logic_1164.all; 
use IEEE.std_logic_unsigned.all; 
use ieee.numeric_std.all;

entity bootloader_dp_32 is
  port (
    CLK:              in std_logic;
    WEA:  in std_logic;
    ENA:  in std_logic;
    MASKA:    in std_logic_vector(3 downto 0);
    ADDRA:         in std_logic_vector(11 downto 2);
    DIA:        in std_logic_vector(31 downto 0);
    DOA:         out std_logic_vector(31 downto 0);
    WEB:  in std_logic;
    ENB:  in std_logic;
    ADDRB:         in std_logic_vector(11 downto 2);
    DIB:        in std_logic_vector(31 downto 0);
    MASKB:    in std_logic_vector(3 downto 0);
    DOB:         out std_logic_vector(31 downto 0)
  );
end entity bootloader_dp_32;

architecture behave of bootloader_dp_32 is

  subtype RAM_WORD is STD_LOGIC_VECTOR (31 downto 0);
  type RAM_TABLE is array (0 to 1023) of RAM_WORD;
 shared variable RAM: RAM_TABLE := RAM_TABLE'(
x"0b0b0b9b",x"af040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b9b",x"99040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fd0608",x"72830609",x"81058205",x"832b2a83",x"ffff0652",x"04000000",x"00000000",x"00000000",x"71fd0608",x"83ffff73",x"83060981",x"05820583",x"2b2b0906",x"7383ffff",x"0b0b0b0b",x"83a70400",x"72098105",x"72057373",x"09060906",x"73097306",x"070a8106",x"53510400",x"00000000",x"00000000",x"72722473",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71737109",x"71068106",x"30720a10",x"0a720a10",x"0a31050a",x"81065151",x"53510400",x"00000000",x"72722673",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"cc040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"720a722b",x"0a535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72729f06",x"0981050b",x"0b0b88af",x"05040000",x"00000000",x"00000000",x"00000000",x"00000000",x"72722aff",x"739f062a",x"0974090a",x"8106ff05",x"06075351",x"04000000",x"00000000",x"00000000",x"71715351",x"020d0406",x"73830609",x"81058205",x"832b0b2b",x"0772fc06",x"0c515104",x"00000000",x"72098105",x"72050970",x"81050906",x"0a810653",x"51040000",x"00000000",x"00000000",x"00000000",x"72098105",x"72050970",x"81050906",x"0a098106",x"53510400",x"00000000",x"00000000",x"00000000",x"71098105",x"52040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72720981",x"05055351",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097206",x"73730906",x"07535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fc0608",x"72830609",x"81058305",x"1010102a",x"81ff0652",x"04000000",x"00000000",x"00000000",x"71fc0608",x"0b0b0b9d",x"ec738306",x"10100508",x"060b0b0b",x"88b20400",x"00000000",x"00000000",x"0b0b0b89",x"80040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"e8040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097081",x"0509060a",x"8106ff05",x"70547106",x"73097274",x"05ff0506",x"07515151",x"04000000",x"72097081",x"0509060a",x"098106ff",x"05705471",x"06730972",x"7405ff05",x"06075151",x"51040000",x"05ff0504",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"810b0b0b",x"0b9eb00c",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71810552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"02840572",x"10100552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"717105ff",x"05715351",x"020d0400",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"81d53f95",x"c53f0400",x"00000000",x"00000000",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101053",x"51047381",x"ff067383",x"06098105",x"83051010",x"102b0772",x"fc060c51",x"51043c04",x"72728072",x"8106ff05",x"09720605",x"71105272",x"0a100a53",x"72ed3851",x"51535104",x"88088c08",x"90087575",x"9cc42d50",x"50880856",x"900c8c0c",x"880c5104",x"88088c08",x"90087575",x"9c892d50",x"50880856",x"900c8c0c",x"880c5104",x"88088c08",x"90088eb3",x"2d900c8c",x"0c880c04",x"ff3d0d0b",x"0b0b9ed4",x"3351709e",x"389ebc08",x"70085252",x"70802e8a",x"3884129e",x"bc0c702d",x"ec39810b",x"0b0b0b9e",x"d434833d",x"0d040480",x"3d0d0b0b",x"0b9f8808",x"802e9738",x"0b0b0b0b",x"800b802e",x"8d380b0b",x"0b9f8851",x"0b0b0bf6",x"873f823d",x"0d0404ff",x"3d0d80c4",x"80808452",x"71087082",x"2a708106",x"51515170",x"f338833d",x"0d04ff3d",x"0d80c480",x"80845271",x"0870812a",x"70810651",x"515170f3",x"38738290",x"0a0c833d",x"0d04fe3d",x"0d747080",x"dc808088",x"0c7081ff",x"06ff8311",x"54515371",x"81268d38",x"80fd518a",x"9a2d72a0",x"32518339",x"72518a9a",x"2d843d0d",x"04ff3d0d",x"028f0533",x"5283ffff",x"0b83d00a",x"0c80fe51",x"8a9a2d71",x"518aba2d",x"833d0d04",x"fe3d0d83",x"d00a0870",x"81ff0652",x"528aba2d",x"71882a51",x"8aba2d80",x"fe518a9a",x"2d9eec33",x"81058706",x"52719eec",x"34843d0d",x"04fe3d0d",x"9ef03370",x"832b8207",x"81fa0652",x"538ae92d",x"8b882d84",x"3d0d04fe",x"3d0d9ef0",x"3370832b",x"810781f9",x"0652538a",x"e92d8b88",x"2d843d0d",x"0482f6ff",x"0b80cc80",x"80880c80",x"0b80cc80",x"80840c9f",x"0b83900a",x"0c04ff3d",x"0d737008",x"515180c8",x"80808470",x"08708480",x"8007720c",x"5252833d",x"0d04ff3d",x"0d80c880",x"80847008",x"70fbffff",x"06720c52",x"52833d0d",x"04a0900b",x"80c0800c",x"9ed80b80",x"c0840c9b",x"902dff3d",x"0d73518b",x"710c9011",x"52988080",x"720c8072",x"0c700883",x"ffff0688",x"0c833d0d",x"04fa3d0d",x"787a7dff",x"1e565658",x"5572ff2e",x"a7388056",x"84527575",x"0c740888",x"180cff12",x"5271f338",x"73841576",x"08720cff",x"15555552",x"72ff2e09",x"8106dd38",x"883d0d04",x"f93d0d80",x"d0808084",x"5783d00a",x"588c9e2d",x"76518cc6",x"2d9ed870",x"88088429",x"98808405",x"71708405",x"530c5656",x"fb8084a1",x"ad750c9e",x"c00b8817",x"0c807078",x"0c770c76",x"087083ff",x"ff065156",x"83ffff78",x"0ca08054",x"88085377",x"5276518c",x"e52d7651",x"8c822d77",x"08557575",x"2e893880",x"c3518a9a",x"2dff39a0",x"84085574",x"fba090ae",x"802e8938",x"80c2518a",x"9a2dff39",x"80d00a70",x"0870ffbf",x"06720c56",x"5689ff2d",x"8cb52dff",x"3d0d9ee4",x"0881119e",x"e40c5183",x"900a7008",x"70feff06",x"720c5252",x"833d0d04",x"fe3d0d9e",x"ec337083",x"2b818007",x"9ef03371",x"81f80607",x"5353538a",x"e92d7481",x"8007518a",x"ba2d8b88",x"2d843d0d",x"04fe3d0d",x"80d08080",x"84538c9e",x"2d85730c",x"80730c72",x"087081ff",x"06745351",x"528c822d",x"71880c84",x"3d0d04fc",x"3d0d7653",x"8bb52d81",x"13338214",x"33718180",x"0a297184",x"80802905",x"83163370",x"82802912",x"84183352",x"7105a080",x"05861885",x"19335952",x"53535456",x"54ff1353",x"72ff2e91",x"38737081",x"05553352",x"71757081",x"055734e9",x"3989518e",x"d02d863d",x"0d04f93d",x"0d795680",x"d0808084",x"578c9e2d",x"81163382",x"17337182",x"80290553",x"5371802e",x"94388516",x"72555372",x"70810554",x"33770cff",x"145473f3",x"38831633",x"84173371",x"82802905",x"56528054",x"73752797",x"38735877",x"770c7316",x"77085353",x"71733481",x"14547474",x"26ed3876",x"518c822d",x"9eec3370",x"832b8180",x"079ef033",x"7181f806",x"07535354",x"8ae92d81",x"84518aba",x"2d74882a",x"518aba2d",x"74518aba",x"2d805473",x"75278f38",x"73167033",x"52528aba",x"2d811454",x"ee398b88",x"2d893d0d",x"04fc3d0d",x"80d08080",x"840b8118",x"54558bb5",x"2d8c9e2d",x"86750c74",x"518c822d",x"8c9e2d82",x"750c7270",x"81055433",x"750c7270",x"81055433",x"750c7270",x"81055433",x"750c81ff",x"54727081",x"05543375",x"0cff1454",x"738025f1",x"3874518c",x"822d8ef9",x"2d880881",x"065271f6",x"38863d0d",x"04fa3d0d",x"785680d0",x"80808454",x"8c9e2d86",x"740c7351",x"8c822d8c",x"9e2d81ad",x"740c8116",x"33821733",x"71828029",x"05831833",x"760c8418",x"33760c85",x"1833760c",x"58528055",x"747727af",x"3874802e",x"88388c9e",x"2d81ad74",x"0c741686",x"1133750c",x"87113375",x"0c527351",x"8c822d8e",x"f92d8808",x"81065271",x"f6388215",x"55ce398c",x"9e2d8474",x"0c73518c",x"822d9eec",x"3370832b",x"8180079e",x"f0337181",x"f8060753",x"53538ae9",x"2d818751",x"8aba2d8b",x"882d883d",x"0d04fc3d",x"0d768111",x"33821233",x"71902b71",x"882b0783",x"14337072",x"07882b84",x"16337107",x"51525356",x"57555288",x"518ed02d",x"81ff518a",x"9a2d80c4",x"80808454",x"73087081",x"2a708106",x"51515271",x"f3387284",x"80800780",x"c4808084",x"0c863d0d",x"04fd3d0d",x"8ef92d88",x"08880881",x"06535371",x"f3389eec",x"3370832b",x"8180079e",x"f0337181",x"f8060753",x"53548ae9",x"2d818351",x"8aba2d72",x"518aba2d",x"8b882d85",x"3d0d04fc",x"3d0d800b",x"9ee40c80",x"709dfc57",x"54547470",x"84055608",x"5271802e",x"8a388113",x"81712b75",x"07555281",x"13538c73",x"27e43873",x"9eec3370",x"832b8180",x"079ef033",x"7181f806",x"07545455",x"538ae92d",x"8181518a",x"ba2d9ec0",x"54935273",x"70810555",x"33518aba",x"2dff1252",x"71ff2e09",x"8106ec38",x"72982a51",x"8aba2d72",x"902a518a",x"ba2d7288",x"2a518aba",x"2d72518a",x"ba2d8051",x"8aba2d8f",x"518aba2d",x"9ec2518a",x"ba2dbd84",x"c0518aba",x"2d8b882d",x"863d0d04",x"fe3d0d80",x"0b9ee40c",x"9eec3370",x"832b8180",x"079ef033",x"7181f806",x"07535353",x"8ae92d81",x"82518aba",x"2d80d080",x"8084528c",x"9e2d81f9",x"0a0b80d0",x"80809c0c",x"71087252",x"538c822d",x"729ef40c",x"72902a51",x"8aba2d9e",x"f408882a",x"518aba2d",x"9ef40851",x"8aba2d8e",x"f92d8808",x"518aba2d",x"8b882d84",x"3d0d0480",x"3d0d810b",x"9ee80c80",x"0b83900a",x"0c85518e",x"d02d823d",x"0d04803d",x"0d800b9e",x"e80c8be9",x"2d86518e",x"d02d823d",x"0d04fd3d",x"0d80d080",x"8084548a",x"518ed02d",x"8c9e2d9e",x"d8745253",x"8cc62d72",x"88088429",x"98808405",x"71708405",x"530c52fb",x"8084a1ad",x"720c9ec0",x"0b88140c",x"73518c82",x"2d89ff2d",x"8cb52dff",x"b23d0d80",x"d23d0856",x"800b9ee8",x"0c800b9e",x"e40c800b",x"df80179e",x"c571902a",x"71565657",x"55577272",x"70810554",x"3473882a",x"53727234",x"73821634",x"75982a52",x"718b1634",x"75902a52",x"718c1634",x"75882a52",x"718d1634",x"758e1634",x"8eb30b80",x"c0800c84",x"80b30b80",x"c4808084",x"0c80c880",x"80a453fb",x"ffff7308",x"70720675",x"0c535480",x"c8808094",x"70087076",x"06720c53",x"53880b80",x"c0808084",x"0c810b90",x"0a0c8be9",x"2dfe8888",x"0b80dc80",x"80840c81",x"f20b80d0",x"0a0c80d0",x"80808470",x"52528c82",x"2d8c9e2d",x"71518c82",x"2d8c9e2d",x"84720c71",x"518c822d",x"76775654",x"80c48080",x"84087081",x"06515271",x"9e389ee8",x"085372ec",x"389ee408",x"5287e872",x"27e23872",x"900a0c72",x"83900a0c",x"9b882d82",x"900a0853",x"74802e81",x"c9387280",x"fe2e0981",x"06818238",x"76802eff",x"bb388055",x"827727ff",x"b33883d0",x"0a085271",x"752e0981",x"06b73888",x"3d337087",x"2a813253",x"5371802e",x"97387287",x"065271ff",x"8f38749e",x"f034749e",x"ec348bb5",x"2dff8139",x"72b80670",x"832a9ef0",x"33555152",x"71732e87",x"388bcf2d",x"feea3981",x"13870652",x"719ef034",x"029d0533",x"52718d26",x"fed63871",x"84299df8",x"0580d13d",x"fde10552",x"70085152",x"712dfec0",x"397280fd",x"2e098106",x"86388154",x"feb23976",x"829f26a5",x"3873802e",x"87388073",x"a0325454",x"7280dc80",x"80880c80",x"d03d7705",x"fde00552",x"72723481",x"1757fe88",x"398055fe",x"83397280",x"fe2e0981",x"06fdf938",x"7457ff0b",x"83d00a0c",x"81775555",x"fdea39ff",x"3d0d9bdd",x"2d735280",x"51979b2d",x"833d0d04",x"83fffff8",x"0d8da004",x"83fffff8",x"0d80c088",x"04880880",x"c0808088",x"0880c080",x"082d5088",x"0c810b90",x"0a0c0480",x"700cfaad",x"95b4da0b",x"81808071",x"710c7180",x"082e8738",x"7011519b",x"bb04519a",x"f72d0000",x"820b80c0",x"8080900c",x"0b0b0b04",x"0083f00a",x"0b800ba0",x"80721208",x"720c8412",x"5271712e",x"ff05f238",x"028c050d",x"9bd00400",x"00000000",x"00000000",x"00000000",x"00fb3d0d",x"77795555",x"80567476",x"25863874",x"30558156",x"73802588",x"38733076",x"81325754",x"80537352",x"745180ca",x"3f880854",x"75802e85",x"38880830",x"5473880c",x"873d0d04",x"fa3d0d78",x"7a575580",x"57747725",x"86387430",x"55815775",x"9f2c5481",x"53757432",x"74315274",x"51943f88",x"08547680",x"2e853888",x"08305473",x"880c883d",x"0d04fc3d",x"0d767853",x"54815380",x"55873971",x"10731054",x"52737226",x"5172802e",x"a7387080",x"2e863871",x"8025e838",x"72802e98",x"38717426",x"89387372",x"31757407",x"56547281",x"2a72812a",x"5353e539",x"73517883",x"38745170",x"880c863d",x"0d04ff3d",x"0d9efc0b",x"fc055271",x"08ff2e8b",x"38710851",x"702dfc12",x"52f13983",x"3d0d0404",x"ebbe3f04",x"00ffffff",x"ff00ffff",x"ffff00ff",x"ffffff00",x"00000a27",x"00000ac4",x"000009ed",x"000007f6",x"00000b2f",x"00000b46",x"000008fd",x"0000099a",x"0000079f",x"00000b5a",x"0000089d",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000f84",x"02010600",x"00000000",x"05b8d800",x"b4041700",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"ffffffff",x"00000000",x"ffffffff",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000");

begin

  process (clk)
  begin
    if rising_edge(clk) then
      if ENA='1' then
        if WEA='1' then
          RAM(conv_integer(ADDRA) ) := DIA;
        end if;
        DOA <= RAM(conv_integer(ADDRA)) ;
      end if;
    end if;
  end process;  

  process (clk)
  begin
    if rising_edge(clk) then
      if ENB='1' then
        if WEB='1' then
          RAM( conv_integer(ADDRB) ) := DIB;
        end if;
        DOB <= RAM(conv_integer(ADDRB)) ;
      end if;
    end if;
  end process;  
end behave;
