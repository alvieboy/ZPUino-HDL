library IEEE;
use IEEE.std_logic_1164.all; 
use IEEE.std_logic_unsigned.all; 
use ieee.numeric_std.all;

entity bootloader_dp_32 is
  port (
    CLK:              in std_logic;
    WEA:  in std_logic;
    ENA:  in std_logic;
    MASKA:    in std_logic_vector(3 downto 0);
    ADDRA:         in std_logic_vector(11 downto 2);
    DIA:        in std_logic_vector(31 downto 0);
    DOA:         out std_logic_vector(31 downto 0);
    WEB:  in std_logic;
    ENB:  in std_logic;
    ADDRB:         in std_logic_vector(11 downto 2);
    DIB:        in std_logic_vector(31 downto 0);
    MASKB:    in std_logic_vector(3 downto 0);
    DOB:         out std_logic_vector(31 downto 0)
  );
end entity bootloader_dp_32;

architecture behave of bootloader_dp_32 is

  subtype RAM_WORD is STD_LOGIC_VECTOR (31 downto 0);
  type RAM_TABLE is array (0 to 1023) of RAM_WORD;
 shared variable RAM: RAM_TABLE := RAM_TABLE'(
x"0b0b0b97",x"8e040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b97",x"af040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fd0608",x"72830609",x"81058205",x"832b2a83",x"ffff0652",x"04000000",x"00000000",x"00000000",x"71fd0608",x"83ffff73",x"83060981",x"05820583",x"2b2b0906",x"7383ffff",x"0b0b0b0b",x"83a70400",x"72098105",x"72057373",x"09060906",x"73097306",x"070a8106",x"53510400",x"00000000",x"00000000",x"72722473",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71737109",x"71068106",x"30720a10",x"0a720a10",x"0a31050a",x"81065151",x"53510400",x"00000000",x"72722673",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"cc040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"720a722b",x"0a535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72729f06",x"0981050b",x"0b0b88af",x"05040000",x"00000000",x"00000000",x"00000000",x"00000000",x"72722aff",x"739f062a",x"0974090a",x"8106ff05",x"06075351",x"04000000",x"00000000",x"00000000",x"71715351",x"020d0406",x"73830609",x"81058205",x"832b0b2b",x"0772fc06",x"0c515104",x"00000000",x"72098105",x"72050970",x"81050906",x"0a810653",x"51040000",x"00000000",x"00000000",x"00000000",x"72098105",x"72050970",x"81050906",x"0a098106",x"53510400",x"00000000",x"00000000",x"00000000",x"71098105",x"52040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72720981",x"05055351",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097206",x"73730906",x"07535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fc0608",x"72830609",x"81058305",x"1010102a",x"81ff0652",x"04000000",x"00000000",x"00000000",x"71fc0608",x"0b0b0b9d",x"cc738306",x"10100508",x"060b0b0b",x"88b20400",x"00000000",x"00000000",x"0b0b0b89",x"80040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"e8040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097081",x"0509060a",x"8106ff05",x"70547106",x"73097274",x"05ff0506",x"07515151",x"04000000",x"72097081",x"0509060a",x"098106ff",x"05705471",x"06730972",x"7405ff05",x"06075151",x"51040000",x"05ff0504",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"810b0b0b",x"0b9e940c",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71810552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"02840572",x"10100552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"717105ff",x"05715351",x"020d0400",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"81dd3f95",x"9a3f0400",x"00000000",x"00000000",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101053",x"51047381",x"ff067383",x"06098105",x"83051010",x"102b0772",x"fc060c51",x"51043c04",x"72728072",x"8106ff05",x"09720605",x"71105272",x"0a100a53",x"72ed3851",x"51535104",x"88088c08",x"90087575",x"98cd2d50",x"50880856",x"900c8c0c",x"880c5104",x"88088c08",x"90087575",x"98892d50",x"50880856",x"900c8c0c",x"880c5104",x"88088c08",x"90088e87",x"2d900c8c",x"0c880c04",x"ff3d0d0b",x"0b0b9ea4",x"335170a6",x"389ea008",x"70085252",x"70802e92",x"3884129e",x"a00c702d",x"9ea00870",x"08525270",x"f038810b",x"0b0b0b9e",x"a434833d",x"0d040480",x"3d0d0b0b",x"0b9ed008",x"802e8e38",x"0b0b0b0b",x"800b802e",x"09810685",x"38823d0d",x"040b0b0b",x"9ed0510b",x"0b0bf5f8",x"3f823d0d",x"0404ff3d",x"0d80c480",x"80845271",x"0870822a",x"70810651",x"515170f3",x"38833d0d",x"04ff3d0d",x"80c48080",x"84527108",x"70812a70",x"81065151",x"5170f338",x"7382900a",x"0c833d0d",x"04fe3d0d",x"747080dc",x"8080880c",x"7081ff06",x"ff831154",x"51537181",x"268d3880",x"fd518aa9",x"2d72a032",x"51833972",x"518aa92d",x"843d0d04",x"803d0d83",x"ffff0b83",x"d00a0c80",x"fe518aa9",x"2d823d0d",x"04ff3d0d",x"83d00a08",x"70882a52",x"528ac92d",x"7181ff06",x"518ac92d",x"80fe518a",x"a92d833d",x"0d0482df",x"c70b80cc",x"8080880c",x"800b80cc",x"8080840c",x"9f0b8390",x"0a0c8e87",x"0ba0800c",x"810b900a",x"0c04ff3d",x"0d737008",x"51518190",x"0a700870",x"820a0772",x"0c525283",x"3d0d04ff",x"3d0d8190",x"0a700870",x"fd0a0672",x"0c525283",x"3d0d04a0",x"900ba080",x"0c9ea80b",x"a0840c97",x"a72dff3d",x"0d73518b",x"710c9011",x"5280dc80",x"80720c80",x"720c7008",x"83ffff06",x"880c833d",x"0d04fa3d",x"0d787a7d",x"ff1e5757",x"585373ff",x"2ea73880",x"56845275",x"730c7208",x"88180cff",x"125271f3",x"38748416",x"7408720c",x"ff165656",x"5273ff2e",x"098106dd",x"38883d0d",x"04f83d0d",x"80d08080",x"845783d0",x"0a598beb",x"2d76518c",x"8e2d9ea8",x"70880810",x"1080dc80",x"84057170",x"8405530c",x"5656fb80",x"84a1ad75",x"0c9e840b",x"88170c80",x"70780c77",x"0c760883",x"ffff0656",x"8fffdf80",x"0b880827",x"8338ff39",x"83ffff79",x"0ca08054",x"88085378",x"5276518c",x"ae2d7651",x"8bd22d78",x"08557476",x"2e893880",x"c3518aa9",x"2dff39a0",x"84085574",x"fbc084b2",x"802e8938",x"80c2518a",x"a92dff39",x"80d00a70",x"0870ffbf",x"06720c56",x"568a8e2d",x"8bff2dff",x"3d0d9eb4",x"0881119e",x"b40c5183",x"900a7008",x"70feff06",x"720c5252",x"833d0d04",x"803d0d8a",x"f82d7281",x"8007518a",x"c92d8b8d",x"2d823d0d",x"04fe3d0d",x"80d08080",x"84538beb",x"2d85730c",x"80730c72",x"087081ff",x"06745351",x"528bd22d",x"71880c84",x"3d0d04fc",x"3d0d7681",x"11338212",x"33718180",x"0a297184",x"80802905",x"83143370",x"82802912",x"84163352",x"7105a080",x"05861685",x"17335752",x"53535557",x"5553ff13",x"5372ff2e",x"91387370",x"81055533",x"52717570",x"81055734",x"e9398951",x"8ea42d86",x"3d0d04f9",x"3d0d7957",x"80d08080",x"84568beb",x"2d811733",x"82183371",x"82802905",x"53537180",x"2e943885",x"17725553",x"72708105",x"5433760c",x"ff145473",x"f3388317",x"33841833",x"71828029",x"05565280",x"54737527",x"97387358",x"77760c73",x"17760853",x"53717334",x"81145474",x"7426ed38",x"75518bd2",x"2d8af82d",x"8184518a",x"c92d7488",x"2a518ac9",x"2d74518a",x"c92d8054",x"7375278f",x"38731770",x"3352528a",x"c92d8114",x"54ee398b",x"8d2d893d",x"0d0404fc",x"3d0d7681",x"11338212",x"3371902b",x"71882b07",x"83143370",x"7207882b",x"84163371",x"07515253",x"57575452",x"88518ea4",x"2d81ff51",x"8aa92d80",x"c4808084",x"53720870",x"812a7081",x"06515152",x"71f33873",x"84808007",x"80c48080",x"840c863d",x"0d04fe3d",x"0d8eb92d",x"88088808",x"81065353",x"71f3388a",x"f82d8183",x"518ac92d",x"72518ac9",x"2d8b8d2d",x"843d0d04",x"fe3d0d80",x"0b9eb40c",x"8af82d81",x"81518ac9",x"2d9e8453",x"8f527270",x"81055433",x"518ac92d",x"ff125271",x"ff2e0981",x"06ec388b",x"8d2d843d",x"0d04fe3d",x"0d800b9e",x"b40c8af8",x"2d818251",x"8ac92d80",x"d0808084",x"528beb2d",x"81f90a0b",x"80d08080",x"9c0c7108",x"7252538b",x"d22d729e",x"bc0c7290",x"2a518ac9",x"2d9ebc08",x"882a518a",x"c92d9ebc",x"08518ac9",x"2d8eb92d",x"8808518a",x"c92d8b8d",x"2d843d0d",x"04803d0d",x"810b9eb8",x"0c800b83",x"900a0c85",x"518ea42d",x"823d0d04",x"803d0d80",x"0b9eb80c",x"8bae2d86",x"518ea42d",x"823d0d04",x"fd3d0d80",x"d0808084",x"548a518e",x"a42d8beb",x"2d9ea874",x"52538c8e",x"2d728808",x"101080dc",x"80840571",x"70840553",x"0c52fb80",x"84a1ad72",x"0c9e840b",x"88140c73",x"518bd22d",x"8a8e2d8b",x"ff2dfc3d",x"0d80d080",x"80847052",x"558bd22d",x"8beb2d8b",x"750c7680",x"d0808094",x"0c80750c",x"a0805477",x"5383d00a",x"5274518c",x"ae2d7451",x"8bd22d8a",x"8e2d8bff",x"2dffab3d",x"0d800b9e",x"b80c800b",x"9eb40c80",x"0b8e870b",x"a0800c57",x"80c48080",x"84558480",x"af750c80",x"c88080a0",x"53fd0a73",x"08707206",x"750c5354",x"80c88080",x"90700870",x"7606720c",x"5353a870",x"99857170",x"8405530c",x"99e2710c",x"539afb0b",x"88120c9c",x"8a0b8c12",x"0c93b60b",x"90120c53",x"880b80c0",x"8080840c",x"900a5381",x"730c8bae",x"2dfe8888",x"0b80dc80",x"80840c81",x"f20b80d0",x"0a0c80d0",x"80808470",x"52528bd2",x"2d8beb2d",x"71518bd2",x"2d767776",x"75933d41",x"415b5b5b",x"83d00a5c",x"78087081",x"06515271",x"9d389eb8",x"085372f0",x"389eb408",x"5287e872",x"27e63872",x"7e0c7283",x"900a0c97",x"9f2d8290",x"0a085379",x"802e81b4",x"387280fe",x"2e098106",x"80f43876",x"802ec138",x"807d7858",x"565a8277",x"27ffb538",x"83ffff7c",x"0c79fe18",x"53537972",x"27983880",x"dc808088",x"72555872",x"15703379",x"0c528113",x"53737326",x"f238ff16",x"75115475",x"05ff0570",x"33743370",x"72882b07",x"7f085351",x"55515271",x"732e0981",x"06feed38",x"74335372",x"8a26fee4",x"38721010",x"9dd80575",x"52700851",x"52712dfe",x"d3397280",x"fd2e0981",x"06863881",x"5bfec539",x"76829f26",x"9e387a80",x"2e873880",x"73a03254",x"5b80d73d",x"7705fde0",x"05527272",x"34811757",x"fea23980",x"5afe9d39",x"7280fe2e",x"098106fe",x"93387957",x"ff7c0c81",x"775c5afe",x"8739ff3d",x"0d97dd2d",x"80528051",x"93ed2d83",x"3d0d048f",x"fffff80d",x"8ce9048f",x"fffff80d",x"a0880488",x"0880c080",x"808808a0",x"80082d50",x"880c810b",x"900a0c04",x"00000000",x"00000000",x"00000000",x"820b80c0",x"8080900c",x"0b0b0b04",x"0083f00a",x"0b800ba0",x"80721208",x"720c8412",x"5271712e",x"ff05f238",x"028c050d",x"97d00400",x"00000000",x"00000000",x"00000000",x"00fb3d0d",x"77795555",x"80567575",x"24ab3880",x"74249d38",x"80537352",x"745180e1",x"3f880854",x"75802e85",x"38880830",x"5473880c",x"873d0d04",x"73307681",x"325754dc",x"39743055",x"81567380",x"25d238ec",x"39fa3d0d",x"787a5755",x"80577675",x"24a43875",x"9f2c5481",x"53757432",x"74315274",x"519b3f88",x"08547680",x"2e853888",x"08305473",x"880c883d",x"0d047430",x"558157d7",x"39fc3d0d",x"76785354",x"81538074",x"73265255",x"72802e98",x"3870802e",x"a9388072",x"24a43871",x"10731075",x"72265354",x"5272ea38",x"73517883",x"38745170",x"880c863d",x"0d047281",x"2a72812a",x"53537280",x"2ee63871",x"7426ef38",x"73723175",x"74077481",x"2a74812a",x"55555654",x"e539fc3d",x"0d767079",x"7b555555",x"558f7227",x"8c387275",x"07830651",x"70802ea7",x"38ff1252",x"71ff2e98",x"38727081",x"05543374",x"70810556",x"34ff1252",x"71ff2e09",x"8106ea38",x"74880c86",x"3d0d0474",x"51727084",x"05540871",x"70840553",x"0c727084",x"05540871",x"70840553",x"0c727084",x"05540871",x"70840553",x"0c727084",x"05540871",x"70840553",x"0cf01252",x"718f26c9",x"38837227",x"95387270",x"84055408",x"71708405",x"530cfc12",x"52718326",x"ed387054",x"ff8339fc",x"3d0d7679",x"71028c05",x"9f053357",x"55535583",x"72278a38",x"74830651",x"70802ea2",x"38ff1252",x"71ff2e93",x"38737370",x"81055534",x"ff125271",x"ff2e0981",x"06ef3874",x"880c863d",x"0d047474",x"882b7507",x"7071902b",x"07515451",x"8f7227a5",x"38727170",x"8405530c",x"72717084",x"05530c72",x"71708405",x"530c7271",x"70840553",x"0cf01252",x"718f26dd",x"38837227",x"90387271",x"70840553",x"0cfc1252",x"718326f2",x"387053ff",x"9039fb3d",x"0d777970",x"72078306",x"53545270",x"93387173",x"73085456",x"54717308",x"2e80c438",x"73755452",x"71337081",x"ff065254",x"70802e9d",x"38723355",x"70752e09",x"81069538",x"81128114",x"71337081",x"ff065456",x"545270e5",x"38723355",x"7381ff06",x"7581ff06",x"71713188",x"0c525287",x"3d0d0471",x"0970f7fb",x"fdff1406",x"70f88482",x"81800651",x"51517097",x"38841484",x"16710854",x"56547175",x"082edc38",x"73755452",x"ff963980",x"0b880c87",x"3d0d04ff",x"3d0d9ec4",x"0bfc0570",x"08525270",x"ff2e9138",x"702dfc12",x"70085252",x"70ff2e09",x"8106f138",x"833d0d04",x"04ebe13f",x"04000000",x"00ffffff",x"ff00ffff",x"ffff00ff",x"ffffff00",x"000008c0",x"000008f2",x"0000089a",x"000007b3",x"00000949",x"00000960",x"00000846",x"00000847",x"0000075f",x"00000974",x"01091700",x"00ffef80",x"055d4a80",x"b8011900",x"00000000",x"00000000",x"00000000",x"00000f4c",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"ffffffff",x"00000000",x"ffffffff",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000");

begin

  process (clk)
  begin
    if rising_edge(clk) then
      if ENA='1' then
        if WEA='1' then
          RAM(conv_integer(ADDRA) ) := DIA;
        end if;
        DOA <= RAM(conv_integer(ADDRA)) ;
      end if;
    end if;
  end process;  

  process (clk)
  begin
    if rising_edge(clk) then
      if ENB='1' then
        if WEB='1' then
          RAM( conv_integer(ADDRB) ) := DIB;
        end if;
        DOB <= RAM(conv_integer(ADDRB)) ;
      end if;
    end if;
  end process;  
end behave;
