library IEEE;
use IEEE.std_logic_1164.all; 
use IEEE.std_logic_unsigned.all; 
use ieee.numeric_std.all;

entity bootloader_dp_32 is
  port (
    CLK:              in std_logic;
    WEA:  in std_logic;
    ENA:  in std_logic;
    MASKA:    in std_logic_vector(3 downto 0);
    ADDRA:         in std_logic_vector(11 downto 2);
    DIA:        in std_logic_vector(31 downto 0);
    DOA:         out std_logic_vector(31 downto 0);
    WEB:  in std_logic;
    ENB:  in std_logic;
    ADDRB:         in std_logic_vector(11 downto 2);
    DIB:        in std_logic_vector(31 downto 0);
    MASKB:    in std_logic_vector(3 downto 0);
    DOB:         out std_logic_vector(31 downto 0)
  );
end entity bootloader_dp_32;

architecture behave of bootloader_dp_32 is

  subtype RAM_WORD is STD_LOGIC_VECTOR (31 downto 0);
  type RAM_TABLE is array (0 to 1023) of RAM_WORD;
 shared variable RAM: RAM_TABLE := RAM_TABLE'(
x"0b0b0b98",x"a0040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b98",x"c1040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fd0608",x"72830609",x"81058205",x"832b2a83",x"ffff0652",x"04000000",x"00000000",x"00000000",x"71fd0608",x"83ffff73",x"83060981",x"05820583",x"2b2b0906",x"7383ffff",x"0b0b0b0b",x"83a70400",x"72098105",x"72057373",x"09060906",x"73097306",x"070a8106",x"53510400",x"00000000",x"00000000",x"72722473",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71737109",x"71068106",x"30720a10",x"0a720a10",x"0a31050a",x"81065151",x"53510400",x"00000000",x"72722673",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"cc040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"720a722b",x"0a535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72729f06",x"0981050b",x"0b0b88af",x"05040000",x"00000000",x"00000000",x"00000000",x"00000000",x"72722aff",x"739f062a",x"0974090a",x"8106ff05",x"06075351",x"04000000",x"00000000",x"00000000",x"71715351",x"020d0406",x"73830609",x"81058205",x"832b0b2b",x"0772fc06",x"0c515104",x"00000000",x"72098105",x"72050970",x"81050906",x"0a810653",x"51040000",x"00000000",x"00000000",x"00000000",x"72098105",x"72050970",x"81050906",x"0a098106",x"53510400",x"00000000",x"00000000",x"00000000",x"71098105",x"52040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72720981",x"05055351",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097206",x"73730906",x"07535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fc0608",x"72830609",x"81058305",x"1010102a",x"81ff0652",x"04000000",x"00000000",x"00000000",x"71fc0608",x"0b0b0b9e",x"dc738306",x"10100508",x"060b0b0b",x"88b20400",x"00000000",x"00000000",x"0b0b0b89",x"80040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"e8040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097081",x"0509060a",x"8106ff05",x"70547106",x"73097274",x"05ff0506",x"07515151",x"04000000",x"72097081",x"0509060a",x"098106ff",x"05705471",x"06730972",x"7405ff05",x"06075151",x"51040000",x"05ff0504",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"810b0b0b",x"0b9fa40c",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71810552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"02840572",x"10100552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"717105ff",x"05715351",x"020d0400",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"81dd3f96",x"aa3f0400",x"00000000",x"00000000",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101053",x"51047381",x"ff067383",x"06098105",x"83051010",x"102b0772",x"fc060c51",x"51043c04",x"72728072",x"8106ff05",x"09720605",x"71105272",x"0a100a53",x"72ed3851",x"51535104",x"88088c08",x"90087575",x"99dd2d50",x"50880856",x"900c8c0c",x"880c5104",x"88088c08",x"90087575",x"99992d50",x"50880856",x"900c8c0c",x"880c5104",x"88088c08",x"90088e80",x"2d900c8c",x"0c880c04",x"ff3d0d0b",x"0b0b9fb4",x"335170a6",x"389fb008",x"70085252",x"70802e92",x"3884129f",x"b00c702d",x"9fb00870",x"08525270",x"f038810b",x"0b0b0b9f",x"b434833d",x"0d040480",x"3d0d0b0b",x"0b9fe008",x"802e8e38",x"0b0b0b0b",x"800b802e",x"09810685",x"38823d0d",x"040b0b0b",x"9fe0510b",x"0b0bf5f8",x"3f823d0d",x"0404ff3d",x"0d80c480",x"80845271",x"0870822a",x"70810651",x"515170f3",x"38833d0d",x"04ff3d0d",x"80c48080",x"84527108",x"70812a70",x"81065151",x"5170f338",x"7382900a",x"0c833d0d",x"04fe3d0d",x"747080dc",x"8080880c",x"7081ff06",x"ff831154",x"51537181",x"268d3880",x"fd518aa9",x"2d72a032",x"51833972",x"518aa92d",x"843d0d04",x"803d0d83",x"ffff0b83",x"d00a0c80",x"fe518aa9",x"2d823d0d",x"04ff3d0d",x"83d00a08",x"70882a52",x"528ac92d",x"7181ff06",x"518ac92d",x"80fe518a",x"a92d833d",x"0d0482f6",x"ff0b80cc",x"8080880c",x"800b80cc",x"8080840c",x"9f0b8390",x"0a0c04ff",x"3d0d7370",x"08515180",x"c8808084",x"70087084",x"80800772",x"0c525283",x"3d0d04ff",x"3d0d80c8",x"80808470",x"0870fbff",x"ff06720c",x"5252833d",x"0d04a090",x"0ba0800c",x"9fb80ba0",x"840c98b9",x"2dff3d0d",x"73518b71",x"0c901152",x"98808072",x"0c80720c",x"700883ff",x"ff06880c",x"833d0d04",x"fa3d0d78",x"7a7dff1e",x"57575853",x"73ff2ea7",x"38805684",x"5275730c",x"72088818",x"0cff1252",x"71f33874",x"84167408",x"720cff16",x"56565273",x"ff2e0981",x"06dd3888",x"3d0d04f8",x"3d0d80d0",x"80808457",x"83d00a59",x"8be32d76",x"518c892d",x"9fb87088",x"08101098",x"80840571",x"70840553",x"0c5656fb",x"8084a1ad",x"750c9f94",x"0b88170c",x"8070780c",x"770c7608",x"83ffff06",x"5683ffdf",x"800b8808",x"278338ff",x"3983ffff",x"790ca080",x"54880853",x"78527651",x"8ca82d76",x"518bc72d",x"78085574",x"762e8938",x"80c3518a",x"a92dff39",x"a0840855",x"74fba090",x"ae802e89",x"3880c251",x"8aa92dff",x"3980d00a",x"700870ff",x"bf06720c",x"56568a8e",x"2d8bfa2d",x"ff3d0d9f",x"c4088111",x"9fc40c51",x"83900a70",x"0870feff",x"06720c52",x"52833d0d",x"04803d0d",x"8af82d72",x"81800751",x"8ac92d8b",x"8d2d823d",x"0d04fe3d",x"0d80d080",x"8084538b",x"e32d8573",x"0c80730c",x"72087081",x"ff067453",x"51528bc7",x"2d71880c",x"843d0d04",x"fc3d0d76",x"81113382",x"12337181",x"800a2971",x"84808029",x"05831433",x"70828029",x"12841633",x"527105a0",x"80058616",x"85173357",x"52535355",x"575553ff",x"135372ff",x"2e913873",x"70810555",x"33527175",x"70810557",x"34e93989",x"518e9d2d",x"863d0d04",x"f93d0d79",x"5780d080",x"8084568b",x"e32d8117",x"33821833",x"71828029",x"05535371",x"802e9438",x"85177255",x"53727081",x"05543376",x"0cff1454",x"73f33883",x"17338418",x"33718280",x"29055652",x"80547375",x"27973873",x"5877760c",x"73177608",x"53537173",x"34811454",x"747426ed",x"3875518b",x"c72d8af8",x"2d818451",x"8ac92d74",x"882a518a",x"c92d7451",x"8ac92d80",x"54737527",x"8f387317",x"70335252",x"8ac92d81",x"1454ee39",x"8b8d2d89",x"3d0d04f9",x"3d0d7956",x"80d08080",x"84558be3",x"2d86750c",x"74518bc7",x"2d8be32d",x"81ad7076",x"0c811733",x"82183371",x"82802905",x"83193378",x"0c841933",x"780c8519",x"33780c59",x"53538054",x"737727b3",x"38725873",x"802e8738",x"8be32d77",x"750c7316",x"86113376",x"0c871133",x"760c5274",x"518bc72d",x"8eb22d88",x"08810652",x"71f63882",x"14547674",x"26d1388b",x"e32d8475",x"0c74518b",x"c72d8af8",x"2d818751",x"8ac92d8b",x"8d2d893d",x"0d04fc3d",x"0d768111",x"33821233",x"71902b71",x"882b0783",x"14337072",x"07882b84",x"16337107",x"51525357",x"57545288",x"518e9d2d",x"81ff518a",x"a92d80c4",x"80808453",x"72087081",x"2a708106",x"51515271",x"f3387384",x"80800780",x"c4808084",x"0c863d0d",x"04fe3d0d",x"8eb22d88",x"08880881",x"06535371",x"f3388af8",x"2d818351",x"8ac92d72",x"518ac92d",x"8b8d2d84",x"3d0d04fe",x"3d0d800b",x"9fc40c8a",x"f82d8181",x"518ac92d",x"9f94538f",x"52727081",x"05543351",x"8ac92dff",x"125271ff",x"2e098106",x"ec388b8d",x"2d843d0d",x"04fe3d0d",x"800b9fc4",x"0c8af82d",x"8182518a",x"c92d80d0",x"80808452",x"8be32d81",x"f90a0b80",x"d080809c",x"0c710872",x"52538bc7",x"2d729fcc",x"0c72902a",x"518ac92d",x"9fcc0888",x"2a518ac9",x"2d9fcc08",x"518ac92d",x"8eb22d88",x"08518ac9",x"2d8b8d2d",x"843d0d04",x"803d0d81",x"0b9fc80c",x"800b8390",x"0a0c8551",x"8e9d2d82",x"3d0d0480",x"3d0d800b",x"9fc80c8b",x"ae2d8651",x"8e9d2d82",x"3d0d04fd",x"3d0d80d0",x"80808454",x"8a518e9d",x"2d8be32d",x"9fb87452",x"538c892d",x"72880810",x"10988084",x"05717084",x"05530c52",x"fb8084a1",x"ad720c9f",x"940b8814",x"0c73518b",x"c72d8a8e",x"2d8bfa2d",x"fc3d0d80",x"d0808084",x"7052558b",x"c72d8be3",x"2d8b750c",x"7680d080",x"80940c80",x"750ca080",x"54775383",x"d00a5274",x"518ca82d",x"74518bc7",x"2d8a8e2d",x"8bfa2dff",x"ab3d0d80",x"0b9fc80c",x"800b9fc4",x"0c800b8e",x"800ba080",x"0c5780c4",x"80808455",x"8480b375",x"0c80c880",x"80a453fb",x"ffff7308",x"70720675",x"0c535480",x"c8808094",x"70087076",x"06720c53",x"53a8709a",x"95717084",x"05530c9a",x"f2710c53",x"9c8b0b88",x"120c9d9a",x"0b8c120c",x"94bc0b90",x"120c5388",x"0b80c080",x"80840c90",x"0a538173",x"0c8bae2d",x"fe88880b",x"80dc8080",x"840c81f2",x"0b80d00a",x"0c80d080",x"80847052",x"528bc72d",x"8be32d71",x"518bc72d",x"8be32d84",x"720c7151",x"8bc72d76",x"77767593",x"3d41415b",x"5b5b83d0",x"0a5c7808",x"70810651",x"52719d38",x"9fc80853",x"72f0389f",x"c4085287",x"e87227e6",x"38727e0c",x"7283900a",x"0c98b12d",x"82900a08",x"5379802e",x"81b43872",x"80fe2e09",x"810680f4",x"3876802e",x"c138807d",x"7858565a",x"827727ff",x"b53883ff",x"ff7c0c79",x"fe185353",x"79722798",x"3880dc80",x"80887255",x"58721570",x"33790c52",x"81135373",x"7326f238",x"ff167511",x"547505ff",x"05703374",x"33707288",x"2b077f08",x"53515551",x"5271732e",x"098106fe",x"ed387433",x"53728a26",x"fee43872",x"10109ee8",x"05755270",x"08515271",x"2dfed339",x"7280fd2e",x"09810686",x"38815bfe",x"c5397682",x"9f269e38",x"7a802e87",x"388073a0",x"32545b80",x"d73d7705",x"fde00552",x"72723481",x"1757fea2",x"39805afe",x"9d397280",x"fe2e0981",x"06fe9338",x"7957ff7c",x"0c81775c",x"5afe8739",x"ff3d0d98",x"ed2d8052",x"805194f3",x"2d833d0d",x"0483ffff",x"f80d8ce3",x"0483ffff",x"f80da088",x"04880880",x"c0808088",x"08a08008",x"2d50880c",x"810b900a",x"0c040000",x"00000000",x"00000000",x"820b80c0",x"8080900c",x"0b0b0b04",x"0083f00a",x"0b800ba0",x"80721208",x"720c8412",x"5271712e",x"ff05f238",x"028c050d",x"98e00400",x"00000000",x"00000000",x"00000000",x"00fb3d0d",x"77795555",x"80567575",x"24ab3880",x"74249d38",x"80537352",x"745180e1",x"3f880854",x"75802e85",x"38880830",x"5473880c",x"873d0d04",x"73307681",x"325754dc",x"39743055",x"81567380",x"25d238ec",x"39fa3d0d",x"787a5755",x"80577675",x"24a43875",x"9f2c5481",x"53757432",x"74315274",x"519b3f88",x"08547680",x"2e853888",x"08305473",x"880c883d",x"0d047430",x"558157d7",x"39fc3d0d",x"76785354",x"81538074",x"73265255",x"72802e98",x"3870802e",x"a9388072",x"24a43871",x"10731075",x"72265354",x"5272ea38",x"73517883",x"38745170",x"880c863d",x"0d047281",x"2a72812a",x"53537280",x"2ee63871",x"7426ef38",x"73723175",x"74077481",x"2a74812a",x"55555654",x"e539fc3d",x"0d767079",x"7b555555",x"558f7227",x"8c387275",x"07830651",x"70802ea7",x"38ff1252",x"71ff2e98",x"38727081",x"05543374",x"70810556",x"34ff1252",x"71ff2e09",x"8106ea38",x"74880c86",x"3d0d0474",x"51727084",x"05540871",x"70840553",x"0c727084",x"05540871",x"70840553",x"0c727084",x"05540871",x"70840553",x"0c727084",x"05540871",x"70840553",x"0cf01252",x"718f26c9",x"38837227",x"95387270",x"84055408",x"71708405",x"530cfc12",x"52718326",x"ed387054",x"ff8339fc",x"3d0d7679",x"71028c05",x"9f053357",x"55535583",x"72278a38",x"74830651",x"70802ea2",x"38ff1252",x"71ff2e93",x"38737370",x"81055534",x"ff125271",x"ff2e0981",x"06ef3874",x"880c863d",x"0d047474",x"882b7507",x"7071902b",x"07515451",x"8f7227a5",x"38727170",x"8405530c",x"72717084",x"05530c72",x"71708405",x"530c7271",x"70840553",x"0cf01252",x"718f26dd",x"38837227",x"90387271",x"70840553",x"0cfc1252",x"718326f2",x"387053ff",x"9039fb3d",x"0d777970",x"72078306",x"53545270",x"93387173",x"73085456",x"54717308",x"2e80c438",x"73755452",x"71337081",x"ff065254",x"70802e9d",x"38723355",x"70752e09",x"81069538",x"81128114",x"71337081",x"ff065456",x"545270e5",x"38723355",x"7381ff06",x"7581ff06",x"71713188",x"0c525287",x"3d0d0471",x"0970f7fb",x"fdff1406",x"70f88482",x"81800651",x"51517097",x"38841484",x"16710854",x"56547175",x"082edc38",x"73755452",x"ff963980",x"0b880c87",x"3d0d04ff",x"3d0d9fd4",x"0bfc0570",x"08525270",x"ff2e9138",x"702dfc12",x"70085252",x"70ff2e09",x"8106f138",x"833d0d04",x"04ead13f",x"04000000",x"00ffffff",x"ff00ffff",x"ffff00ff",x"ffffff00",x"00000947",x"00000979",x"00000921",x"000007ac",x"000009d0",x"000009e7",x"0000083f",x"000008ce",x"00000758",x"000009fb",x"01090600",x"007fef80",x"05b8d800",x"b4041700",x"00000000",x"00000000",x"00000000",x"00000fdc",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"ffffffff",x"00000000",x"ffffffff",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000");

begin

  process (clk)
  begin
    if rising_edge(clk) then
      if ENA='1' then
        if WEA='1' then
          RAM(conv_integer(ADDRA) ) := DIA;
        end if;
        DOA <= RAM(conv_integer(ADDRA)) ;
      end if;
    end if;
  end process;  

  process (clk)
  begin
    if rising_edge(clk) then
      if ENB='1' then
        if WEB='1' then
          RAM( conv_integer(ADDRB) ) := DIB;
        end if;
        DOB <= RAM(conv_integer(ADDRB)) ;
      end if;
    end if;
  end process;  
end behave;
