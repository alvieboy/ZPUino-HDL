---------------------------------------------------------------------
--	Filename:	gh_sincos_rom_12.vhd
--			
--	Description:
--		Sin Cos look up table 12 bit 
--
--	Copyright (c) 2008 by George Huber 
--		an OpenCores.org Project
--		free to use, but see documentation for conditions 
--
--	Revision 	History:
--	Revision 	Date      	Author   	Comment
--	-------- 	----------	---------	-----------
--	1.0      	10/26/08  	h LeFevre	Initial revision
--	
------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

entity gh_sincos_rom_12 is
	port (
		CLK : in std_logic;
		ADD : in std_logic_vector(11 downto 0);
		sin : out std_logic_vector(11 downto 0);
		cos : out std_logic_vector(11 downto 0)
		);
end entity;

architecture a of gh_sincos_rom_12 is

	type rom_mem is array (0 to 4095) of std_logic_vector (11 downto 0);
	constant isin : rom_mem :=(  
    x"000", x"003", x"006", x"009", x"00d", x"010", x"013", x"016", 
    x"019", x"01c", x"01f", x"023", x"026", x"029", x"02c", x"02f", 
    x"032", x"035", x"039", x"03c", x"03f", x"042", x"045", x"048", 
    x"04b", x"04e", x"052", x"055", x"058", x"05b", x"05e", x"061", 
    x"064", x"068", x"06b", x"06e", x"071", x"074", x"077", x"07a", 
    x"07e", x"081", x"084", x"087", x"08a", x"08d", x"090", x"093", 
    x"097", x"09a", x"09d", x"0a0", x"0a3", x"0a6", x"0a9", x"0ac", 
    x"0b0", x"0b3", x"0b6", x"0b9", x"0bc", x"0bf", x"0c2", x"0c6", 
    x"0c9", x"0cc", x"0cf", x"0d2", x"0d5", x"0d8", x"0db", x"0df", 
    x"0e2", x"0e5", x"0e8", x"0eb", x"0ee", x"0f1", x"0f4", x"0f7", 
    x"0fb", x"0fe", x"101", x"104", x"107", x"10a", x"10d", x"110", 
    x"113", x"117", x"11a", x"11d", x"120", x"123", x"126", x"129", 
    x"12c", x"12f", x"133", x"136", x"139", x"13c", x"13f", x"142", 
    x"145", x"148", x"14b", x"14e", x"152", x"155", x"158", x"15b", 
    x"15e", x"161", x"164", x"167", x"16a", x"16d", x"171", x"174", 
    x"177", x"17a", x"17d", x"180", x"183", x"186", x"189", x"18c", 
    x"18f", x"192", x"196", x"199", x"19c", x"19f", x"1a2", x"1a5", 
    x"1a8", x"1ab", x"1ae", x"1b1", x"1b4", x"1b7", x"1ba", x"1bd", 
    x"1c1", x"1c4", x"1c7", x"1ca", x"1cd", x"1d0", x"1d3", x"1d6", 
    x"1d9", x"1dc", x"1df", x"1e2", x"1e5", x"1e8", x"1eb", x"1ee", 
    x"1f1", x"1f4", x"1f7", x"1fb", x"1fe", x"201", x"204", x"207", 
    x"20a", x"20d", x"210", x"213", x"216", x"219", x"21c", x"21f", 
    x"222", x"225", x"228", x"22b", x"22e", x"231", x"234", x"237", 
    x"23a", x"23d", x"240", x"243", x"246", x"249", x"24c", x"24f", 
    x"252", x"255", x"258", x"25b", x"25e", x"261", x"264", x"267", 
    x"26a", x"26d", x"270", x"273", x"276", x"279", x"27c", x"27f", 
    x"282", x"285", x"288", x"28b", x"28e", x"291", x"294", x"297", 
    x"29a", x"29d", x"2a0", x"2a3", x"2a6", x"2a9", x"2ac", x"2af", 
    x"2b2", x"2b5", x"2b8", x"2ba", x"2bd", x"2c0", x"2c3", x"2c6", 
    x"2c9", x"2cc", x"2cf", x"2d2", x"2d5", x"2d8", x"2db", x"2de", 
    x"2e1", x"2e4", x"2e7", x"2e9", x"2ec", x"2ef", x"2f2", x"2f5", 
    x"2f8", x"2fb", x"2fe", x"301", x"304", x"307", x"30a", x"30c", 
    x"30f", x"312", x"315", x"318", x"31b", x"31e", x"321", x"324", 
    x"327", x"329", x"32c", x"32f", x"332", x"335", x"338", x"33b", 
    x"33e", x"340", x"343", x"346", x"349", x"34c", x"34f", x"352", 
    x"354", x"357", x"35a", x"35d", x"360", x"363", x"366", x"368", 
    x"36b", x"36e", x"371", x"374", x"377", x"379", x"37c", x"37f", 
    x"382", x"385", x"387", x"38a", x"38d", x"390", x"393", x"396", 
    x"398", x"39b", x"39e", x"3a1", x"3a4", x"3a6", x"3a9", x"3ac", 
    x"3af", x"3b2", x"3b4", x"3b7", x"3ba", x"3bd", x"3bf", x"3c2", 
    x"3c5", x"3c8", x"3ca", x"3cd", x"3d0", x"3d3", x"3d6", x"3d8", 
    x"3db", x"3de", x"3e1", x"3e3", x"3e6", x"3e9", x"3eb", x"3ee", 
    x"3f1", x"3f4", x"3f6", x"3f9", x"3fc", x"3ff", x"401", x"404", 
    x"407", x"409", x"40c", x"40f", x"412", x"414", x"417", x"41a", 
    x"41c", x"41f", x"422", x"424", x"427", x"42a", x"42c", x"42f", 
    x"432", x"435", x"437", x"43a", x"43d", x"43f", x"442", x"444", 
    x"447", x"44a", x"44c", x"44f", x"452", x"454", x"457", x"45a", 
    x"45c", x"45f", x"462", x"464", x"467", x"469", x"46c", x"46f", 
    x"471", x"474", x"476", x"479", x"47c", x"47e", x"481", x"483", 
    x"486", x"489", x"48b", x"48e", x"490", x"493", x"496", x"498", 
    x"49b", x"49d", x"4a0", x"4a2", x"4a5", x"4a7", x"4aa", x"4ad", 
    x"4af", x"4b2", x"4b4", x"4b7", x"4b9", x"4bc", x"4be", x"4c1", 
    x"4c3", x"4c6", x"4c8", x"4cb", x"4cd", x"4d0", x"4d2", x"4d5", 
    x"4d7", x"4da", x"4dc", x"4df", x"4e1", x"4e4", x"4e6", x"4e9", 
    x"4eb", x"4ee", x"4f0", x"4f3", x"4f5", x"4f8", x"4fa", x"4fd", 
    x"4ff", x"502", x"504", x"506", x"509", x"50b", x"50e", x"510", 
    x"513", x"515", x"517", x"51a", x"51c", x"51f", x"521", x"524", 
    x"526", x"528", x"52b", x"52d", x"530", x"532", x"534", x"537", 
    x"539", x"53b", x"53e", x"540", x"543", x"545", x"547", x"54a", 
    x"54c", x"54e", x"551", x"553", x"555", x"558", x"55a", x"55c", 
    x"55f", x"561", x"563", x"566", x"568", x"56a", x"56d", x"56f", 
    x"571", x"573", x"576", x"578", x"57a", x"57d", x"57f", x"581", 
    x"583", x"586", x"588", x"58a", x"58d", x"58f", x"591", x"593", 
    x"596", x"598", x"59a", x"59c", x"59f", x"5a1", x"5a3", x"5a5", 
    x"5a7", x"5aa", x"5ac", x"5ae", x"5b0", x"5b3", x"5b5", x"5b7", 
    x"5b9", x"5bb", x"5bd", x"5c0", x"5c2", x"5c4", x"5c6", x"5c8", 
    x"5cb", x"5cd", x"5cf", x"5d1", x"5d3", x"5d5", x"5d7", x"5da", 
    x"5dc", x"5de", x"5e0", x"5e2", x"5e4", x"5e6", x"5e9", x"5eb", 
    x"5ed", x"5ef", x"5f1", x"5f3", x"5f5", x"5f7", x"5f9", x"5fb", 
    x"5fd", x"600", x"602", x"604", x"606", x"608", x"60a", x"60c", 
    x"60e", x"610", x"612", x"614", x"616", x"618", x"61a", x"61c", 
    x"61e", x"620", x"622", x"624", x"626", x"628", x"62a", x"62c", 
    x"62e", x"630", x"632", x"634", x"636", x"638", x"63a", x"63c", 
    x"63e", x"640", x"642", x"644", x"646", x"648", x"64a", x"64c", 
    x"64e", x"650", x"652", x"654", x"655", x"657", x"659", x"65b", 
    x"65d", x"65f", x"661", x"663", x"665", x"667", x"668", x"66a", 
    x"66c", x"66e", x"670", x"672", x"674", x"675", x"677", x"679", 
    x"67b", x"67d", x"67f", x"681", x"682", x"684", x"686", x"688", 
    x"68a", x"68b", x"68d", x"68f", x"691", x"693", x"694", x"696", 
    x"698", x"69a", x"69b", x"69d", x"69f", x"6a1", x"6a3", x"6a4", 
    x"6a6", x"6a8", x"6a9", x"6ab", x"6ad", x"6af", x"6b0", x"6b2", 
    x"6b4", x"6b6", x"6b7", x"6b9", x"6bb", x"6bc", x"6be", x"6c0", 
    x"6c1", x"6c3", x"6c5", x"6c6", x"6c8", x"6ca", x"6cb", x"6cd", 
    x"6cf", x"6d0", x"6d2", x"6d4", x"6d5", x"6d7", x"6d9", x"6da", 
    x"6dc", x"6dd", x"6df", x"6e1", x"6e2", x"6e4", x"6e5", x"6e7", 
    x"6e9", x"6ea", x"6ec", x"6ed", x"6ef", x"6f0", x"6f2", x"6f4", 
    x"6f5", x"6f7", x"6f8", x"6fa", x"6fb", x"6fd", x"6fe", x"700", 
    x"701", x"703", x"704", x"706", x"707", x"709", x"70a", x"70c", 
    x"70d", x"70f", x"710", x"712", x"713", x"715", x"716", x"718", 
    x"719", x"71a", x"71c", x"71d", x"71f", x"720", x"722", x"723", 
    x"724", x"726", x"727", x"729", x"72a", x"72b", x"72d", x"72e", 
    x"730", x"731", x"732", x"734", x"735", x"736", x"738", x"739", 
    x"73a", x"73c", x"73d", x"73e", x"740", x"741", x"742", x"744", 
    x"745", x"746", x"748", x"749", x"74a", x"74c", x"74d", x"74e", 
    x"74f", x"751", x"752", x"753", x"754", x"756", x"757", x"758", 
    x"759", x"75b", x"75c", x"75d", x"75e", x"760", x"761", x"762", 
    x"763", x"764", x"766", x"767", x"768", x"769", x"76a", x"76b", 
    x"76d", x"76e", x"76f", x"770", x"771", x"772", x"774", x"775", 
    x"776", x"777", x"778", x"779", x"77a", x"77b", x"77d", x"77e", 
    x"77f", x"780", x"781", x"782", x"783", x"784", x"785", x"786", 
    x"787", x"788", x"789", x"78a", x"78c", x"78d", x"78e", x"78f", 
    x"790", x"791", x"792", x"793", x"794", x"795", x"796", x"797", 
    x"798", x"799", x"79a", x"79b", x"79c", x"79d", x"79e", x"79e", 
    x"79f", x"7a0", x"7a1", x"7a2", x"7a3", x"7a4", x"7a5", x"7a6", 
    x"7a7", x"7a8", x"7a9", x"7aa", x"7aa", x"7ab", x"7ac", x"7ad", 
    x"7ae", x"7af", x"7b0", x"7b1", x"7b1", x"7b2", x"7b3", x"7b4", 
    x"7b5", x"7b6", x"7b7", x"7b7", x"7b8", x"7b9", x"7ba", x"7bb", 
    x"7bb", x"7bc", x"7bd", x"7be", x"7bf", x"7bf", x"7c0", x"7c1", 
    x"7c2", x"7c2", x"7c3", x"7c4", x"7c5", x"7c5", x"7c6", x"7c7", 
    x"7c8", x"7c8", x"7c9", x"7ca", x"7ca", x"7cb", x"7cc", x"7cd", 
    x"7cd", x"7ce", x"7cf", x"7cf", x"7d0", x"7d1", x"7d1", x"7d2", 
    x"7d3", x"7d3", x"7d4", x"7d5", x"7d5", x"7d6", x"7d6", x"7d7", 
    x"7d8", x"7d8", x"7d9", x"7d9", x"7da", x"7db", x"7db", x"7dc", 
    x"7dc", x"7dd", x"7de", x"7de", x"7df", x"7df", x"7e0", x"7e0", 
    x"7e1", x"7e1", x"7e2", x"7e2", x"7e3", x"7e3", x"7e4", x"7e5", 
    x"7e5", x"7e6", x"7e6", x"7e6", x"7e7", x"7e7", x"7e8", x"7e8", 
    x"7e9", x"7e9", x"7ea", x"7ea", x"7eb", x"7eb", x"7ec", x"7ec", 
    x"7ec", x"7ed", x"7ed", x"7ee", x"7ee", x"7ee", x"7ef", x"7ef", 
    x"7f0", x"7f0", x"7f0", x"7f1", x"7f1", x"7f1", x"7f2", x"7f2", 
    x"7f3", x"7f3", x"7f3", x"7f4", x"7f4", x"7f4", x"7f5", x"7f5", 
    x"7f5", x"7f5", x"7f6", x"7f6", x"7f6", x"7f7", x"7f7", x"7f7", 
    x"7f7", x"7f8", x"7f8", x"7f8", x"7f8", x"7f9", x"7f9", x"7f9", 
    x"7f9", x"7fa", x"7fa", x"7fa", x"7fa", x"7fb", x"7fb", x"7fb", 
    x"7fb", x"7fb", x"7fc", x"7fc", x"7fc", x"7fc", x"7fc", x"7fc", 
    x"7fd", x"7fd", x"7fd", x"7fd", x"7fd", x"7fd", x"7fd", x"7fd", 
    x"7fe", x"7fe", x"7fe", x"7fe", x"7fe", x"7fe", x"7fe", x"7fe", 
    x"7fe", x"7fe", x"7ff", x"7ff", x"7ff", x"7ff", x"7ff", x"7ff", 
    x"7ff", x"7ff", x"7ff", x"7ff", x"7ff", x"7ff", x"7ff", x"7ff", 
    x"7ff", x"7ff", x"7ff", x"7ff", x"7ff", x"7ff", x"7ff", x"7ff", 
    x"7ff", x"7ff", x"7ff", x"7ff", x"7ff", x"7ff", x"7ff", x"7fe", 
    x"7fe", x"7fe", x"7fe", x"7fe", x"7fe", x"7fe", x"7fe", x"7fe", 
    x"7fe", x"7fd", x"7fd", x"7fd", x"7fd", x"7fd", x"7fd", x"7fd", 
    x"7fd", x"7fc", x"7fc", x"7fc", x"7fc", x"7fc", x"7fc", x"7fb", 
    x"7fb", x"7fb", x"7fb", x"7fb", x"7fa", x"7fa", x"7fa", x"7fa", 
    x"7f9", x"7f9", x"7f9", x"7f9", x"7f8", x"7f8", x"7f8", x"7f8", 
    x"7f7", x"7f7", x"7f7", x"7f7", x"7f6", x"7f6", x"7f6", x"7f5", 
    x"7f5", x"7f5", x"7f5", x"7f4", x"7f4", x"7f4", x"7f3", x"7f3", 
    x"7f3", x"7f2", x"7f2", x"7f1", x"7f1", x"7f1", x"7f0", x"7f0", 
    x"7f0", x"7ef", x"7ef", x"7ee", x"7ee", x"7ee", x"7ed", x"7ed", 
    x"7ec", x"7ec", x"7ec", x"7eb", x"7eb", x"7ea", x"7ea", x"7e9", 
    x"7e9", x"7e8", x"7e8", x"7e7", x"7e7", x"7e6", x"7e6", x"7e6", 
    x"7e5", x"7e5", x"7e4", x"7e3", x"7e3", x"7e2", x"7e2", x"7e1", 
    x"7e1", x"7e0", x"7e0", x"7df", x"7df", x"7de", x"7de", x"7dd", 
    x"7dc", x"7dc", x"7db", x"7db", x"7da", x"7d9", x"7d9", x"7d8", 
    x"7d8", x"7d7", x"7d6", x"7d6", x"7d5", x"7d5", x"7d4", x"7d3", 
    x"7d3", x"7d2", x"7d1", x"7d1", x"7d0", x"7cf", x"7cf", x"7ce", 
    x"7cd", x"7cd", x"7cc", x"7cb", x"7ca", x"7ca", x"7c9", x"7c8", 
    x"7c8", x"7c7", x"7c6", x"7c5", x"7c5", x"7c4", x"7c3", x"7c2", 
    x"7c2", x"7c1", x"7c0", x"7bf", x"7bf", x"7be", x"7bd", x"7bc", 
    x"7bb", x"7bb", x"7ba", x"7b9", x"7b8", x"7b7", x"7b7", x"7b6", 
    x"7b5", x"7b4", x"7b3", x"7b2", x"7b1", x"7b1", x"7b0", x"7af", 
    x"7ae", x"7ad", x"7ac", x"7ab", x"7aa", x"7aa", x"7a9", x"7a8", 
    x"7a7", x"7a6", x"7a5", x"7a4", x"7a3", x"7a2", x"7a1", x"7a0", 
    x"79f", x"79e", x"79e", x"79d", x"79c", x"79b", x"79a", x"799", 
    x"798", x"797", x"796", x"795", x"794", x"793", x"792", x"791", 
    x"790", x"78f", x"78e", x"78d", x"78c", x"78a", x"789", x"788", 
    x"787", x"786", x"785", x"784", x"783", x"782", x"781", x"780", 
    x"77f", x"77e", x"77d", x"77b", x"77a", x"779", x"778", x"777", 
    x"776", x"775", x"774", x"772", x"771", x"770", x"76f", x"76e", 
    x"76d", x"76b", x"76a", x"769", x"768", x"767", x"766", x"764", 
    x"763", x"762", x"761", x"760", x"75e", x"75d", x"75c", x"75b", 
    x"759", x"758", x"757", x"756", x"754", x"753", x"752", x"751", 
    x"74f", x"74e", x"74d", x"74c", x"74a", x"749", x"748", x"746", 
    x"745", x"744", x"742", x"741", x"740", x"73e", x"73d", x"73c", 
    x"73a", x"739", x"738", x"736", x"735", x"734", x"732", x"731", 
    x"730", x"72e", x"72d", x"72b", x"72a", x"729", x"727", x"726", 
    x"724", x"723", x"722", x"720", x"71f", x"71d", x"71c", x"71a", 
    x"719", x"718", x"716", x"715", x"713", x"712", x"710", x"70f", 
    x"70d", x"70c", x"70a", x"709", x"707", x"706", x"704", x"703", 
    x"701", x"700", x"6fe", x"6fd", x"6fb", x"6fa", x"6f8", x"6f7", 
    x"6f5", x"6f4", x"6f2", x"6f0", x"6ef", x"6ed", x"6ec", x"6ea", 
    x"6e9", x"6e7", x"6e5", x"6e4", x"6e2", x"6e1", x"6df", x"6dd", 
    x"6dc", x"6da", x"6d9", x"6d7", x"6d5", x"6d4", x"6d2", x"6d0", 
    x"6cf", x"6cd", x"6cb", x"6ca", x"6c8", x"6c6", x"6c5", x"6c3", 
    x"6c1", x"6c0", x"6be", x"6bc", x"6bb", x"6b9", x"6b7", x"6b6", 
    x"6b4", x"6b2", x"6b0", x"6af", x"6ad", x"6ab", x"6a9", x"6a8", 
    x"6a6", x"6a4", x"6a3", x"6a1", x"69f", x"69d", x"69b", x"69a", 
    x"698", x"696", x"694", x"693", x"691", x"68f", x"68d", x"68b", 
    x"68a", x"688", x"686", x"684", x"682", x"681", x"67f", x"67d", 
    x"67b", x"679", x"677", x"675", x"674", x"672", x"670", x"66e", 
    x"66c", x"66a", x"668", x"667", x"665", x"663", x"661", x"65f", 
    x"65d", x"65b", x"659", x"657", x"655", x"654", x"652", x"650", 
    x"64e", x"64c", x"64a", x"648", x"646", x"644", x"642", x"640", 
    x"63e", x"63c", x"63a", x"638", x"636", x"634", x"632", x"630", 
    x"62e", x"62c", x"62a", x"628", x"626", x"624", x"622", x"620", 
    x"61e", x"61c", x"61a", x"618", x"616", x"614", x"612", x"610", 
    x"60e", x"60c", x"60a", x"608", x"606", x"604", x"602", x"600", 
    x"5fd", x"5fb", x"5f9", x"5f7", x"5f5", x"5f3", x"5f1", x"5ef", 
    x"5ed", x"5eb", x"5e9", x"5e6", x"5e4", x"5e2", x"5e0", x"5de", 
    x"5dc", x"5da", x"5d7", x"5d5", x"5d3", x"5d1", x"5cf", x"5cd", 
    x"5cb", x"5c8", x"5c6", x"5c4", x"5c2", x"5c0", x"5bd", x"5bb", 
    x"5b9", x"5b7", x"5b5", x"5b3", x"5b0", x"5ae", x"5ac", x"5aa", 
    x"5a7", x"5a5", x"5a3", x"5a1", x"59f", x"59c", x"59a", x"598", 
    x"596", x"593", x"591", x"58f", x"58d", x"58a", x"588", x"586", 
    x"583", x"581", x"57f", x"57d", x"57a", x"578", x"576", x"573", 
    x"571", x"56f", x"56d", x"56a", x"568", x"566", x"563", x"561", 
    x"55f", x"55c", x"55a", x"558", x"555", x"553", x"551", x"54e", 
    x"54c", x"54a", x"547", x"545", x"543", x"540", x"53e", x"53b", 
    x"539", x"537", x"534", x"532", x"530", x"52d", x"52b", x"528", 
    x"526", x"524", x"521", x"51f", x"51c", x"51a", x"517", x"515", 
    x"513", x"510", x"50e", x"50b", x"509", x"506", x"504", x"502", 
    x"4ff", x"4fd", x"4fa", x"4f8", x"4f5", x"4f3", x"4f0", x"4ee", 
    x"4eb", x"4e9", x"4e6", x"4e4", x"4e1", x"4df", x"4dc", x"4da", 
    x"4d7", x"4d5", x"4d2", x"4d0", x"4cd", x"4cb", x"4c8", x"4c6", 
    x"4c3", x"4c1", x"4be", x"4bc", x"4b9", x"4b7", x"4b4", x"4b2", 
    x"4af", x"4ad", x"4aa", x"4a7", x"4a5", x"4a2", x"4a0", x"49d", 
    x"49b", x"498", x"496", x"493", x"490", x"48e", x"48b", x"489", 
    x"486", x"483", x"481", x"47e", x"47c", x"479", x"476", x"474", 
    x"471", x"46f", x"46c", x"469", x"467", x"464", x"462", x"45f", 
    x"45c", x"45a", x"457", x"454", x"452", x"44f", x"44c", x"44a", 
    x"447", x"444", x"442", x"43f", x"43d", x"43a", x"437", x"435", 
    x"432", x"42f", x"42c", x"42a", x"427", x"424", x"422", x"41f", 
    x"41c", x"41a", x"417", x"414", x"412", x"40f", x"40c", x"409", 
    x"407", x"404", x"401", x"3ff", x"3fc", x"3f9", x"3f6", x"3f4", 
    x"3f1", x"3ee", x"3eb", x"3e9", x"3e6", x"3e3", x"3e1", x"3de", 
    x"3db", x"3d8", x"3d6", x"3d3", x"3d0", x"3cd", x"3ca", x"3c8", 
    x"3c5", x"3c2", x"3bf", x"3bd", x"3ba", x"3b7", x"3b4", x"3b2", 
    x"3af", x"3ac", x"3a9", x"3a6", x"3a4", x"3a1", x"39e", x"39b", 
    x"398", x"396", x"393", x"390", x"38d", x"38a", x"387", x"385", 
    x"382", x"37f", x"37c", x"379", x"377", x"374", x"371", x"36e", 
    x"36b", x"368", x"366", x"363", x"360", x"35d", x"35a", x"357", 
    x"354", x"352", x"34f", x"34c", x"349", x"346", x"343", x"340", 
    x"33e", x"33b", x"338", x"335", x"332", x"32f", x"32c", x"329", 
    x"327", x"324", x"321", x"31e", x"31b", x"318", x"315", x"312", 
    x"30f", x"30c", x"30a", x"307", x"304", x"301", x"2fe", x"2fb", 
    x"2f8", x"2f5", x"2f2", x"2ef", x"2ec", x"2e9", x"2e7", x"2e4", 
    x"2e1", x"2de", x"2db", x"2d8", x"2d5", x"2d2", x"2cf", x"2cc", 
    x"2c9", x"2c6", x"2c3", x"2c0", x"2bd", x"2ba", x"2b8", x"2b5", 
    x"2b2", x"2af", x"2ac", x"2a9", x"2a6", x"2a3", x"2a0", x"29d", 
    x"29a", x"297", x"294", x"291", x"28e", x"28b", x"288", x"285", 
    x"282", x"27f", x"27c", x"279", x"276", x"273", x"270", x"26d", 
    x"26a", x"267", x"264", x"261", x"25e", x"25b", x"258", x"255", 
    x"252", x"24f", x"24c", x"249", x"246", x"243", x"240", x"23d", 
    x"23a", x"237", x"234", x"231", x"22e", x"22b", x"228", x"225", 
    x"222", x"21f", x"21c", x"219", x"216", x"213", x"210", x"20d", 
    x"20a", x"207", x"204", x"201", x"1fe", x"1fb", x"1f7", x"1f4", 
    x"1f1", x"1ee", x"1eb", x"1e8", x"1e5", x"1e2", x"1df", x"1dc", 
    x"1d9", x"1d6", x"1d3", x"1d0", x"1cd", x"1ca", x"1c7", x"1c4", 
    x"1c1", x"1bd", x"1ba", x"1b7", x"1b4", x"1b1", x"1ae", x"1ab", 
    x"1a8", x"1a5", x"1a2", x"19f", x"19c", x"199", x"196", x"192", 
    x"18f", x"18c", x"189", x"186", x"183", x"180", x"17d", x"17a", 
    x"177", x"174", x"171", x"16d", x"16a", x"167", x"164", x"161", 
    x"15e", x"15b", x"158", x"155", x"152", x"14e", x"14b", x"148", 
    x"145", x"142", x"13f", x"13c", x"139", x"136", x"133", x"12f", 
    x"12c", x"129", x"126", x"123", x"120", x"11d", x"11a", x"117", 
    x"113", x"110", x"10d", x"10a", x"107", x"104", x"101", x"0fe", 
    x"0fb", x"0f7", x"0f4", x"0f1", x"0ee", x"0eb", x"0e8", x"0e5", 
    x"0e2", x"0df", x"0db", x"0d8", x"0d5", x"0d2", x"0cf", x"0cc", 
    x"0c9", x"0c6", x"0c2", x"0bf", x"0bc", x"0b9", x"0b6", x"0b3", 
    x"0b0", x"0ac", x"0a9", x"0a6", x"0a3", x"0a0", x"09d", x"09a", 
    x"097", x"093", x"090", x"08d", x"08a", x"087", x"084", x"081", 
    x"07e", x"07a", x"077", x"074", x"071", x"06e", x"06b", x"068", 
    x"064", x"061", x"05e", x"05b", x"058", x"055", x"052", x"04e", 
    x"04b", x"048", x"045", x"042", x"03f", x"03c", x"039", x"035", 
    x"032", x"02f", x"02c", x"029", x"026", x"023", x"01f", x"01c", 
    x"019", x"016", x"013", x"010", x"00d", x"009", x"006", x"003", 
    x"000", x"ffd", x"ffa", x"ff7", x"ff3", x"ff0", x"fed", x"fea", 
    x"fe7", x"fe4", x"fe1", x"fdd", x"fda", x"fd7", x"fd4", x"fd1", 
    x"fce", x"fcb", x"fc7", x"fc4", x"fc1", x"fbe", x"fbb", x"fb8", 
    x"fb5", x"fb2", x"fae", x"fab", x"fa8", x"fa5", x"fa2", x"f9f", 
    x"f9c", x"f98", x"f95", x"f92", x"f8f", x"f8c", x"f89", x"f86", 
    x"f82", x"f7f", x"f7c", x"f79", x"f76", x"f73", x"f70", x"f6d", 
    x"f69", x"f66", x"f63", x"f60", x"f5d", x"f5a", x"f57", x"f54", 
    x"f50", x"f4d", x"f4a", x"f47", x"f44", x"f41", x"f3e", x"f3a", 
    x"f37", x"f34", x"f31", x"f2e", x"f2b", x"f28", x"f25", x"f21", 
    x"f1e", x"f1b", x"f18", x"f15", x"f12", x"f0f", x"f0c", x"f09", 
    x"f05", x"f02", x"eff", x"efc", x"ef9", x"ef6", x"ef3", x"ef0", 
    x"eed", x"ee9", x"ee6", x"ee3", x"ee0", x"edd", x"eda", x"ed7", 
    x"ed4", x"ed1", x"ecd", x"eca", x"ec7", x"ec4", x"ec1", x"ebe", 
    x"ebb", x"eb8", x"eb5", x"eb2", x"eae", x"eab", x"ea8", x"ea5", 
    x"ea2", x"e9f", x"e9c", x"e99", x"e96", x"e93", x"e8f", x"e8c", 
    x"e89", x"e86", x"e83", x"e80", x"e7d", x"e7a", x"e77", x"e74", 
    x"e71", x"e6e", x"e6a", x"e67", x"e64", x"e61", x"e5e", x"e5b", 
    x"e58", x"e55", x"e52", x"e4f", x"e4c", x"e49", x"e46", x"e43", 
    x"e3f", x"e3c", x"e39", x"e36", x"e33", x"e30", x"e2d", x"e2a", 
    x"e27", x"e24", x"e21", x"e1e", x"e1b", x"e18", x"e15", x"e12", 
    x"e0f", x"e0c", x"e09", x"e05", x"e02", x"dff", x"dfc", x"df9", 
    x"df6", x"df3", x"df0", x"ded", x"dea", x"de7", x"de4", x"de1", 
    x"dde", x"ddb", x"dd8", x"dd5", x"dd2", x"dcf", x"dcc", x"dc9", 
    x"dc6", x"dc3", x"dc0", x"dbd", x"dba", x"db7", x"db4", x"db1", 
    x"dae", x"dab", x"da8", x"da5", x"da2", x"d9f", x"d9c", x"d99", 
    x"d96", x"d93", x"d90", x"d8d", x"d8a", x"d87", x"d84", x"d81", 
    x"d7e", x"d7b", x"d78", x"d75", x"d72", x"d6f", x"d6c", x"d69", 
    x"d66", x"d63", x"d60", x"d5d", x"d5a", x"d57", x"d54", x"d51", 
    x"d4e", x"d4b", x"d48", x"d46", x"d43", x"d40", x"d3d", x"d3a", 
    x"d37", x"d34", x"d31", x"d2e", x"d2b", x"d28", x"d25", x"d22", 
    x"d1f", x"d1c", x"d19", x"d17", x"d14", x"d11", x"d0e", x"d0b", 
    x"d08", x"d05", x"d02", x"cff", x"cfc", x"cf9", x"cf6", x"cf4", 
    x"cf1", x"cee", x"ceb", x"ce8", x"ce5", x"ce2", x"cdf", x"cdc", 
    x"cd9", x"cd7", x"cd4", x"cd1", x"cce", x"ccb", x"cc8", x"cc5", 
    x"cc2", x"cc0", x"cbd", x"cba", x"cb7", x"cb4", x"cb1", x"cae", 
    x"cac", x"ca9", x"ca6", x"ca3", x"ca0", x"c9d", x"c9a", x"c98", 
    x"c95", x"c92", x"c8f", x"c8c", x"c89", x"c87", x"c84", x"c81", 
    x"c7e", x"c7b", x"c79", x"c76", x"c73", x"c70", x"c6d", x"c6a", 
    x"c68", x"c65", x"c62", x"c5f", x"c5c", x"c5a", x"c57", x"c54", 
    x"c51", x"c4e", x"c4c", x"c49", x"c46", x"c43", x"c41", x"c3e", 
    x"c3b", x"c38", x"c36", x"c33", x"c30", x"c2d", x"c2a", x"c28", 
    x"c25", x"c22", x"c1f", x"c1d", x"c1a", x"c17", x"c15", x"c12", 
    x"c0f", x"c0c", x"c0a", x"c07", x"c04", x"c01", x"bff", x"bfc", 
    x"bf9", x"bf7", x"bf4", x"bf1", x"bee", x"bec", x"be9", x"be6", 
    x"be4", x"be1", x"bde", x"bdc", x"bd9", x"bd6", x"bd4", x"bd1", 
    x"bce", x"bcb", x"bc9", x"bc6", x"bc3", x"bc1", x"bbe", x"bbc", 
    x"bb9", x"bb6", x"bb4", x"bb1", x"bae", x"bac", x"ba9", x"ba6", 
    x"ba4", x"ba1", x"b9e", x"b9c", x"b99", x"b97", x"b94", x"b91", 
    x"b8f", x"b8c", x"b8a", x"b87", x"b84", x"b82", x"b7f", x"b7d", 
    x"b7a", x"b77", x"b75", x"b72", x"b70", x"b6d", x"b6a", x"b68", 
    x"b65", x"b63", x"b60", x"b5e", x"b5b", x"b59", x"b56", x"b53", 
    x"b51", x"b4e", x"b4c", x"b49", x"b47", x"b44", x"b42", x"b3f", 
    x"b3d", x"b3a", x"b38", x"b35", x"b33", x"b30", x"b2e", x"b2b", 
    x"b29", x"b26", x"b24", x"b21", x"b1f", x"b1c", x"b1a", x"b17", 
    x"b15", x"b12", x"b10", x"b0d", x"b0b", x"b08", x"b06", x"b03", 
    x"b01", x"afe", x"afc", x"afa", x"af7", x"af5", x"af2", x"af0", 
    x"aed", x"aeb", x"ae9", x"ae6", x"ae4", x"ae1", x"adf", x"adc", 
    x"ada", x"ad8", x"ad5", x"ad3", x"ad0", x"ace", x"acc", x"ac9", 
    x"ac7", x"ac5", x"ac2", x"ac0", x"abd", x"abb", x"ab9", x"ab6", 
    x"ab4", x"ab2", x"aaf", x"aad", x"aab", x"aa8", x"aa6", x"aa4", 
    x"aa1", x"a9f", x"a9d", x"a9a", x"a98", x"a96", x"a93", x"a91", 
    x"a8f", x"a8d", x"a8a", x"a88", x"a86", x"a83", x"a81", x"a7f", 
    x"a7d", x"a7a", x"a78", x"a76", x"a73", x"a71", x"a6f", x"a6d", 
    x"a6a", x"a68", x"a66", x"a64", x"a61", x"a5f", x"a5d", x"a5b", 
    x"a59", x"a56", x"a54", x"a52", x"a50", x"a4d", x"a4b", x"a49", 
    x"a47", x"a45", x"a43", x"a40", x"a3e", x"a3c", x"a3a", x"a38", 
    x"a35", x"a33", x"a31", x"a2f", x"a2d", x"a2b", x"a29", x"a26", 
    x"a24", x"a22", x"a20", x"a1e", x"a1c", x"a1a", x"a17", x"a15", 
    x"a13", x"a11", x"a0f", x"a0d", x"a0b", x"a09", x"a07", x"a05", 
    x"a03", x"a00", x"9fe", x"9fc", x"9fa", x"9f8", x"9f6", x"9f4", 
    x"9f2", x"9f0", x"9ee", x"9ec", x"9ea", x"9e8", x"9e6", x"9e4", 
    x"9e2", x"9e0", x"9de", x"9dc", x"9da", x"9d8", x"9d6", x"9d4", 
    x"9d2", x"9d0", x"9ce", x"9cc", x"9ca", x"9c8", x"9c6", x"9c4", 
    x"9c2", x"9c0", x"9be", x"9bc", x"9ba", x"9b8", x"9b6", x"9b4", 
    x"9b2", x"9b0", x"9ae", x"9ac", x"9ab", x"9a9", x"9a7", x"9a5", 
    x"9a3", x"9a1", x"99f", x"99d", x"99b", x"999", x"998", x"996", 
    x"994", x"992", x"990", x"98e", x"98c", x"98b", x"989", x"987", 
    x"985", x"983", x"981", x"97f", x"97e", x"97c", x"97a", x"978", 
    x"976", x"975", x"973", x"971", x"96f", x"96d", x"96c", x"96a", 
    x"968", x"966", x"965", x"963", x"961", x"95f", x"95d", x"95c", 
    x"95a", x"958", x"957", x"955", x"953", x"951", x"950", x"94e", 
    x"94c", x"94a", x"949", x"947", x"945", x"944", x"942", x"940", 
    x"93f", x"93d", x"93b", x"93a", x"938", x"936", x"935", x"933", 
    x"931", x"930", x"92e", x"92c", x"92b", x"929", x"927", x"926", 
    x"924", x"923", x"921", x"91f", x"91e", x"91c", x"91b", x"919", 
    x"917", x"916", x"914", x"913", x"911", x"910", x"90e", x"90c", 
    x"90b", x"909", x"908", x"906", x"905", x"903", x"902", x"900", 
    x"8ff", x"8fd", x"8fc", x"8fa", x"8f9", x"8f7", x"8f6", x"8f4", 
    x"8f3", x"8f1", x"8f0", x"8ee", x"8ed", x"8eb", x"8ea", x"8e8", 
    x"8e7", x"8e6", x"8e4", x"8e3", x"8e1", x"8e0", x"8de", x"8dd", 
    x"8dc", x"8da", x"8d9", x"8d7", x"8d6", x"8d5", x"8d3", x"8d2", 
    x"8d0", x"8cf", x"8ce", x"8cc", x"8cb", x"8ca", x"8c8", x"8c7", 
    x"8c6", x"8c4", x"8c3", x"8c2", x"8c0", x"8bf", x"8be", x"8bc", 
    x"8bb", x"8ba", x"8b8", x"8b7", x"8b6", x"8b4", x"8b3", x"8b2", 
    x"8b1", x"8af", x"8ae", x"8ad", x"8ac", x"8aa", x"8a9", x"8a8", 
    x"8a7", x"8a5", x"8a4", x"8a3", x"8a2", x"8a0", x"89f", x"89e", 
    x"89d", x"89c", x"89a", x"899", x"898", x"897", x"896", x"895", 
    x"893", x"892", x"891", x"890", x"88f", x"88e", x"88c", x"88b", 
    x"88a", x"889", x"888", x"887", x"886", x"885", x"883", x"882", 
    x"881", x"880", x"87f", x"87e", x"87d", x"87c", x"87b", x"87a", 
    x"879", x"878", x"877", x"876", x"874", x"873", x"872", x"871", 
    x"870", x"86f", x"86e", x"86d", x"86c", x"86b", x"86a", x"869", 
    x"868", x"867", x"866", x"865", x"864", x"863", x"862", x"862", 
    x"861", x"860", x"85f", x"85e", x"85d", x"85c", x"85b", x"85a", 
    x"859", x"858", x"857", x"856", x"856", x"855", x"854", x"853", 
    x"852", x"851", x"850", x"84f", x"84f", x"84e", x"84d", x"84c", 
    x"84b", x"84a", x"849", x"849", x"848", x"847", x"846", x"845", 
    x"845", x"844", x"843", x"842", x"841", x"841", x"840", x"83f", 
    x"83e", x"83e", x"83d", x"83c", x"83b", x"83b", x"83a", x"839", 
    x"838", x"838", x"837", x"836", x"836", x"835", x"834", x"833", 
    x"833", x"832", x"831", x"831", x"830", x"82f", x"82f", x"82e", 
    x"82d", x"82d", x"82c", x"82b", x"82b", x"82a", x"82a", x"829", 
    x"828", x"828", x"827", x"827", x"826", x"825", x"825", x"824", 
    x"824", x"823", x"822", x"822", x"821", x"821", x"820", x"820", 
    x"81f", x"81f", x"81e", x"81e", x"81d", x"81d", x"81c", x"81b", 
    x"81b", x"81a", x"81a", x"81a", x"819", x"819", x"818", x"818", 
    x"817", x"817", x"816", x"816", x"815", x"815", x"814", x"814", 
    x"814", x"813", x"813", x"812", x"812", x"812", x"811", x"811", 
    x"810", x"810", x"810", x"80f", x"80f", x"80f", x"80e", x"80e", 
    x"80d", x"80d", x"80d", x"80c", x"80c", x"80c", x"80b", x"80b", 
    x"80b", x"80b", x"80a", x"80a", x"80a", x"809", x"809", x"809", 
    x"809", x"808", x"808", x"808", x"808", x"807", x"807", x"807", 
    x"807", x"806", x"806", x"806", x"806", x"805", x"805", x"805", 
    x"805", x"805", x"804", x"804", x"804", x"804", x"804", x"804", 
    x"803", x"803", x"803", x"803", x"803", x"803", x"803", x"803", 
    x"802", x"802", x"802", x"802", x"802", x"802", x"802", x"802", 
    x"802", x"802", x"801", x"801", x"801", x"801", x"801", x"801", 
    x"801", x"801", x"801", x"801", x"801", x"801", x"801", x"801", 
    x"801", x"801", x"801", x"801", x"801", x"801", x"801", x"801", 
    x"801", x"801", x"801", x"801", x"801", x"801", x"801", x"802", 
    x"802", x"802", x"802", x"802", x"802", x"802", x"802", x"802", 
    x"802", x"803", x"803", x"803", x"803", x"803", x"803", x"803", 
    x"803", x"804", x"804", x"804", x"804", x"804", x"804", x"805", 
    x"805", x"805", x"805", x"805", x"806", x"806", x"806", x"806", 
    x"807", x"807", x"807", x"807", x"808", x"808", x"808", x"808", 
    x"809", x"809", x"809", x"809", x"80a", x"80a", x"80a", x"80b", 
    x"80b", x"80b", x"80b", x"80c", x"80c", x"80c", x"80d", x"80d", 
    x"80d", x"80e", x"80e", x"80f", x"80f", x"80f", x"810", x"810", 
    x"810", x"811", x"811", x"812", x"812", x"812", x"813", x"813", 
    x"814", x"814", x"814", x"815", x"815", x"816", x"816", x"817", 
    x"817", x"818", x"818", x"819", x"819", x"81a", x"81a", x"81a", 
    x"81b", x"81b", x"81c", x"81d", x"81d", x"81e", x"81e", x"81f", 
    x"81f", x"820", x"820", x"821", x"821", x"822", x"822", x"823", 
    x"824", x"824", x"825", x"825", x"826", x"827", x"827", x"828", 
    x"828", x"829", x"82a", x"82a", x"82b", x"82b", x"82c", x"82d", 
    x"82d", x"82e", x"82f", x"82f", x"830", x"831", x"831", x"832", 
    x"833", x"833", x"834", x"835", x"836", x"836", x"837", x"838", 
    x"838", x"839", x"83a", x"83b", x"83b", x"83c", x"83d", x"83e", 
    x"83e", x"83f", x"840", x"841", x"841", x"842", x"843", x"844", 
    x"845", x"845", x"846", x"847", x"848", x"849", x"849", x"84a", 
    x"84b", x"84c", x"84d", x"84e", x"84f", x"84f", x"850", x"851", 
    x"852", x"853", x"854", x"855", x"856", x"856", x"857", x"858", 
    x"859", x"85a", x"85b", x"85c", x"85d", x"85e", x"85f", x"860", 
    x"861", x"862", x"862", x"863", x"864", x"865", x"866", x"867", 
    x"868", x"869", x"86a", x"86b", x"86c", x"86d", x"86e", x"86f", 
    x"870", x"871", x"872", x"873", x"874", x"876", x"877", x"878", 
    x"879", x"87a", x"87b", x"87c", x"87d", x"87e", x"87f", x"880", 
    x"881", x"882", x"883", x"885", x"886", x"887", x"888", x"889", 
    x"88a", x"88b", x"88c", x"88e", x"88f", x"890", x"891", x"892", 
    x"893", x"895", x"896", x"897", x"898", x"899", x"89a", x"89c", 
    x"89d", x"89e", x"89f", x"8a0", x"8a2", x"8a3", x"8a4", x"8a5", 
    x"8a7", x"8a8", x"8a9", x"8aa", x"8ac", x"8ad", x"8ae", x"8af", 
    x"8b1", x"8b2", x"8b3", x"8b4", x"8b6", x"8b7", x"8b8", x"8ba", 
    x"8bb", x"8bc", x"8be", x"8bf", x"8c0", x"8c2", x"8c3", x"8c4", 
    x"8c6", x"8c7", x"8c8", x"8ca", x"8cb", x"8cc", x"8ce", x"8cf", 
    x"8d0", x"8d2", x"8d3", x"8d5", x"8d6", x"8d7", x"8d9", x"8da", 
    x"8dc", x"8dd", x"8de", x"8e0", x"8e1", x"8e3", x"8e4", x"8e6", 
    x"8e7", x"8e8", x"8ea", x"8eb", x"8ed", x"8ee", x"8f0", x"8f1", 
    x"8f3", x"8f4", x"8f6", x"8f7", x"8f9", x"8fa", x"8fc", x"8fd", 
    x"8ff", x"900", x"902", x"903", x"905", x"906", x"908", x"909", 
    x"90b", x"90c", x"90e", x"910", x"911", x"913", x"914", x"916", 
    x"917", x"919", x"91b", x"91c", x"91e", x"91f", x"921", x"923", 
    x"924", x"926", x"927", x"929", x"92b", x"92c", x"92e", x"930", 
    x"931", x"933", x"935", x"936", x"938", x"93a", x"93b", x"93d", 
    x"93f", x"940", x"942", x"944", x"945", x"947", x"949", x"94a", 
    x"94c", x"94e", x"950", x"951", x"953", x"955", x"957", x"958", 
    x"95a", x"95c", x"95d", x"95f", x"961", x"963", x"965", x"966", 
    x"968", x"96a", x"96c", x"96d", x"96f", x"971", x"973", x"975", 
    x"976", x"978", x"97a", x"97c", x"97e", x"97f", x"981", x"983", 
    x"985", x"987", x"989", x"98b", x"98c", x"98e", x"990", x"992", 
    x"994", x"996", x"998", x"999", x"99b", x"99d", x"99f", x"9a1", 
    x"9a3", x"9a5", x"9a7", x"9a9", x"9ab", x"9ac", x"9ae", x"9b0", 
    x"9b2", x"9b4", x"9b6", x"9b8", x"9ba", x"9bc", x"9be", x"9c0", 
    x"9c2", x"9c4", x"9c6", x"9c8", x"9ca", x"9cc", x"9ce", x"9d0", 
    x"9d2", x"9d4", x"9d6", x"9d8", x"9da", x"9dc", x"9de", x"9e0", 
    x"9e2", x"9e4", x"9e6", x"9e8", x"9ea", x"9ec", x"9ee", x"9f0", 
    x"9f2", x"9f4", x"9f6", x"9f8", x"9fa", x"9fc", x"9fe", x"a00", 
    x"a03", x"a05", x"a07", x"a09", x"a0b", x"a0d", x"a0f", x"a11", 
    x"a13", x"a15", x"a17", x"a1a", x"a1c", x"a1e", x"a20", x"a22", 
    x"a24", x"a26", x"a29", x"a2b", x"a2d", x"a2f", x"a31", x"a33", 
    x"a35", x"a38", x"a3a", x"a3c", x"a3e", x"a40", x"a43", x"a45", 
    x"a47", x"a49", x"a4b", x"a4d", x"a50", x"a52", x"a54", x"a56", 
    x"a59", x"a5b", x"a5d", x"a5f", x"a61", x"a64", x"a66", x"a68", 
    x"a6a", x"a6d", x"a6f", x"a71", x"a73", x"a76", x"a78", x"a7a", 
    x"a7d", x"a7f", x"a81", x"a83", x"a86", x"a88", x"a8a", x"a8d", 
    x"a8f", x"a91", x"a93", x"a96", x"a98", x"a9a", x"a9d", x"a9f", 
    x"aa1", x"aa4", x"aa6", x"aa8", x"aab", x"aad", x"aaf", x"ab2", 
    x"ab4", x"ab6", x"ab9", x"abb", x"abd", x"ac0", x"ac2", x"ac5", 
    x"ac7", x"ac9", x"acc", x"ace", x"ad0", x"ad3", x"ad5", x"ad8", 
    x"ada", x"adc", x"adf", x"ae1", x"ae4", x"ae6", x"ae9", x"aeb", 
    x"aed", x"af0", x"af2", x"af5", x"af7", x"afa", x"afc", x"afe", 
    x"b01", x"b03", x"b06", x"b08", x"b0b", x"b0d", x"b10", x"b12", 
    x"b15", x"b17", x"b1a", x"b1c", x"b1f", x"b21", x"b24", x"b26", 
    x"b29", x"b2b", x"b2e", x"b30", x"b33", x"b35", x"b38", x"b3a", 
    x"b3d", x"b3f", x"b42", x"b44", x"b47", x"b49", x"b4c", x"b4e", 
    x"b51", x"b53", x"b56", x"b59", x"b5b", x"b5e", x"b60", x"b63", 
    x"b65", x"b68", x"b6a", x"b6d", x"b70", x"b72", x"b75", x"b77", 
    x"b7a", x"b7d", x"b7f", x"b82", x"b84", x"b87", x"b8a", x"b8c", 
    x"b8f", x"b91", x"b94", x"b97", x"b99", x"b9c", x"b9e", x"ba1", 
    x"ba4", x"ba6", x"ba9", x"bac", x"bae", x"bb1", x"bb4", x"bb6", 
    x"bb9", x"bbc", x"bbe", x"bc1", x"bc3", x"bc6", x"bc9", x"bcb", 
    x"bce", x"bd1", x"bd4", x"bd6", x"bd9", x"bdc", x"bde", x"be1", 
    x"be4", x"be6", x"be9", x"bec", x"bee", x"bf1", x"bf4", x"bf7", 
    x"bf9", x"bfc", x"bff", x"c01", x"c04", x"c07", x"c0a", x"c0c", 
    x"c0f", x"c12", x"c15", x"c17", x"c1a", x"c1d", x"c1f", x"c22", 
    x"c25", x"c28", x"c2a", x"c2d", x"c30", x"c33", x"c36", x"c38", 
    x"c3b", x"c3e", x"c41", x"c43", x"c46", x"c49", x"c4c", x"c4e", 
    x"c51", x"c54", x"c57", x"c5a", x"c5c", x"c5f", x"c62", x"c65", 
    x"c68", x"c6a", x"c6d", x"c70", x"c73", x"c76", x"c79", x"c7b", 
    x"c7e", x"c81", x"c84", x"c87", x"c89", x"c8c", x"c8f", x"c92", 
    x"c95", x"c98", x"c9a", x"c9d", x"ca0", x"ca3", x"ca6", x"ca9", 
    x"cac", x"cae", x"cb1", x"cb4", x"cb7", x"cba", x"cbd", x"cc0", 
    x"cc2", x"cc5", x"cc8", x"ccb", x"cce", x"cd1", x"cd4", x"cd7", 
    x"cd9", x"cdc", x"cdf", x"ce2", x"ce5", x"ce8", x"ceb", x"cee", 
    x"cf1", x"cf4", x"cf6", x"cf9", x"cfc", x"cff", x"d02", x"d05", 
    x"d08", x"d0b", x"d0e", x"d11", x"d14", x"d17", x"d19", x"d1c", 
    x"d1f", x"d22", x"d25", x"d28", x"d2b", x"d2e", x"d31", x"d34", 
    x"d37", x"d3a", x"d3d", x"d40", x"d43", x"d46", x"d48", x"d4b", 
    x"d4e", x"d51", x"d54", x"d57", x"d5a", x"d5d", x"d60", x"d63", 
    x"d66", x"d69", x"d6c", x"d6f", x"d72", x"d75", x"d78", x"d7b", 
    x"d7e", x"d81", x"d84", x"d87", x"d8a", x"d8d", x"d90", x"d93", 
    x"d96", x"d99", x"d9c", x"d9f", x"da2", x"da5", x"da8", x"dab", 
    x"dae", x"db1", x"db4", x"db7", x"dba", x"dbd", x"dc0", x"dc3", 
    x"dc6", x"dc9", x"dcc", x"dcf", x"dd2", x"dd5", x"dd8", x"ddb", 
    x"dde", x"de1", x"de4", x"de7", x"dea", x"ded", x"df0", x"df3", 
    x"df6", x"df9", x"dfc", x"dff", x"e02", x"e05", x"e09", x"e0c", 
    x"e0f", x"e12", x"e15", x"e18", x"e1b", x"e1e", x"e21", x"e24", 
    x"e27", x"e2a", x"e2d", x"e30", x"e33", x"e36", x"e39", x"e3c", 
    x"e3f", x"e43", x"e46", x"e49", x"e4c", x"e4f", x"e52", x"e55", 
    x"e58", x"e5b", x"e5e", x"e61", x"e64", x"e67", x"e6a", x"e6e", 
    x"e71", x"e74", x"e77", x"e7a", x"e7d", x"e80", x"e83", x"e86", 
    x"e89", x"e8c", x"e8f", x"e93", x"e96", x"e99", x"e9c", x"e9f", 
    x"ea2", x"ea5", x"ea8", x"eab", x"eae", x"eb2", x"eb5", x"eb8", 
    x"ebb", x"ebe", x"ec1", x"ec4", x"ec7", x"eca", x"ecd", x"ed1", 
    x"ed4", x"ed7", x"eda", x"edd", x"ee0", x"ee3", x"ee6", x"ee9", 
    x"eed", x"ef0", x"ef3", x"ef6", x"ef9", x"efc", x"eff", x"f02", 
    x"f05", x"f09", x"f0c", x"f0f", x"f12", x"f15", x"f18", x"f1b", 
    x"f1e", x"f21", x"f25", x"f28", x"f2b", x"f2e", x"f31", x"f34", 
    x"f37", x"f3a", x"f3e", x"f41", x"f44", x"f47", x"f4a", x"f4d", 
    x"f50", x"f54", x"f57", x"f5a", x"f5d", x"f60", x"f63", x"f66", 
    x"f69", x"f6d", x"f70", x"f73", x"f76", x"f79", x"f7c", x"f7f", 
    x"f82", x"f86", x"f89", x"f8c", x"f8f", x"f92", x"f95", x"f98", 
    x"f9c", x"f9f", x"fa2", x"fa5", x"fa8", x"fab", x"fae", x"fb2", 
    x"fb5", x"fb8", x"fbb", x"fbe", x"fc1", x"fc4", x"fc7", x"fcb", 
    x"fce", x"fd1", x"fd4", x"fd7", x"fda", x"fdd", x"fe1", x"fe4", 
    x"fe7", x"fea", x"fed", x"ff0", x"ff3", x"ff7", x"ffa", x"ffd");

	constant icos : rom_mem :=( 
    x"7ff", x"7ff", x"7ff", x"7ff", x"7ff", x"7ff", x"7ff", x"7ff", 
    x"7ff", x"7ff", x"7ff", x"7ff", x"7ff", x"7ff", x"7ff", x"7fe", 
    x"7fe", x"7fe", x"7fe", x"7fe", x"7fe", x"7fe", x"7fe", x"7fe", 
    x"7fe", x"7fd", x"7fd", x"7fd", x"7fd", x"7fd", x"7fd", x"7fd", 
    x"7fd", x"7fc", x"7fc", x"7fc", x"7fc", x"7fc", x"7fc", x"7fb", 
    x"7fb", x"7fb", x"7fb", x"7fb", x"7fa", x"7fa", x"7fa", x"7fa", 
    x"7f9", x"7f9", x"7f9", x"7f9", x"7f8", x"7f8", x"7f8", x"7f8", 
    x"7f7", x"7f7", x"7f7", x"7f7", x"7f6", x"7f6", x"7f6", x"7f5", 
    x"7f5", x"7f5", x"7f5", x"7f4", x"7f4", x"7f4", x"7f3", x"7f3", 
    x"7f3", x"7f2", x"7f2", x"7f1", x"7f1", x"7f1", x"7f0", x"7f0", 
    x"7f0", x"7ef", x"7ef", x"7ee", x"7ee", x"7ee", x"7ed", x"7ed", 
    x"7ec", x"7ec", x"7ec", x"7eb", x"7eb", x"7ea", x"7ea", x"7e9", 
    x"7e9", x"7e8", x"7e8", x"7e7", x"7e7", x"7e6", x"7e6", x"7e6", 
    x"7e5", x"7e5", x"7e4", x"7e3", x"7e3", x"7e2", x"7e2", x"7e1", 
    x"7e1", x"7e0", x"7e0", x"7df", x"7df", x"7de", x"7de", x"7dd", 
    x"7dc", x"7dc", x"7db", x"7db", x"7da", x"7d9", x"7d9", x"7d8", 
    x"7d8", x"7d7", x"7d6", x"7d6", x"7d5", x"7d5", x"7d4", x"7d3", 
    x"7d3", x"7d2", x"7d1", x"7d1", x"7d0", x"7cf", x"7cf", x"7ce", 
    x"7cd", x"7cd", x"7cc", x"7cb", x"7ca", x"7ca", x"7c9", x"7c8", 
    x"7c8", x"7c7", x"7c6", x"7c5", x"7c5", x"7c4", x"7c3", x"7c2", 
    x"7c2", x"7c1", x"7c0", x"7bf", x"7bf", x"7be", x"7bd", x"7bc", 
    x"7bb", x"7bb", x"7ba", x"7b9", x"7b8", x"7b7", x"7b7", x"7b6", 
    x"7b5", x"7b4", x"7b3", x"7b2", x"7b1", x"7b1", x"7b0", x"7af", 
    x"7ae", x"7ad", x"7ac", x"7ab", x"7aa", x"7aa", x"7a9", x"7a8", 
    x"7a7", x"7a6", x"7a5", x"7a4", x"7a3", x"7a2", x"7a1", x"7a0", 
    x"79f", x"79e", x"79e", x"79d", x"79c", x"79b", x"79a", x"799", 
    x"798", x"797", x"796", x"795", x"794", x"793", x"792", x"791", 
    x"790", x"78f", x"78e", x"78d", x"78c", x"78a", x"789", x"788", 
    x"787", x"786", x"785", x"784", x"783", x"782", x"781", x"780", 
    x"77f", x"77e", x"77d", x"77b", x"77a", x"779", x"778", x"777", 
    x"776", x"775", x"774", x"772", x"771", x"770", x"76f", x"76e", 
    x"76d", x"76b", x"76a", x"769", x"768", x"767", x"766", x"764", 
    x"763", x"762", x"761", x"760", x"75e", x"75d", x"75c", x"75b", 
    x"759", x"758", x"757", x"756", x"754", x"753", x"752", x"751", 
    x"74f", x"74e", x"74d", x"74c", x"74a", x"749", x"748", x"746", 
    x"745", x"744", x"742", x"741", x"740", x"73e", x"73d", x"73c", 
    x"73a", x"739", x"738", x"736", x"735", x"734", x"732", x"731", 
    x"730", x"72e", x"72d", x"72b", x"72a", x"729", x"727", x"726", 
    x"724", x"723", x"722", x"720", x"71f", x"71d", x"71c", x"71a", 
    x"719", x"718", x"716", x"715", x"713", x"712", x"710", x"70f", 
    x"70d", x"70c", x"70a", x"709", x"707", x"706", x"704", x"703", 
    x"701", x"700", x"6fe", x"6fd", x"6fb", x"6fa", x"6f8", x"6f7", 
    x"6f5", x"6f4", x"6f2", x"6f0", x"6ef", x"6ed", x"6ec", x"6ea", 
    x"6e9", x"6e7", x"6e5", x"6e4", x"6e2", x"6e1", x"6df", x"6dd", 
    x"6dc", x"6da", x"6d9", x"6d7", x"6d5", x"6d4", x"6d2", x"6d0", 
    x"6cf", x"6cd", x"6cb", x"6ca", x"6c8", x"6c6", x"6c5", x"6c3", 
    x"6c1", x"6c0", x"6be", x"6bc", x"6bb", x"6b9", x"6b7", x"6b6", 
    x"6b4", x"6b2", x"6b0", x"6af", x"6ad", x"6ab", x"6a9", x"6a8", 
    x"6a6", x"6a4", x"6a3", x"6a1", x"69f", x"69d", x"69b", x"69a", 
    x"698", x"696", x"694", x"693", x"691", x"68f", x"68d", x"68b", 
    x"68a", x"688", x"686", x"684", x"682", x"681", x"67f", x"67d", 
    x"67b", x"679", x"677", x"675", x"674", x"672", x"670", x"66e", 
    x"66c", x"66a", x"668", x"667", x"665", x"663", x"661", x"65f", 
    x"65d", x"65b", x"659", x"657", x"655", x"654", x"652", x"650", 
    x"64e", x"64c", x"64a", x"648", x"646", x"644", x"642", x"640", 
    x"63e", x"63c", x"63a", x"638", x"636", x"634", x"632", x"630", 
    x"62e", x"62c", x"62a", x"628", x"626", x"624", x"622", x"620", 
    x"61e", x"61c", x"61a", x"618", x"616", x"614", x"612", x"610", 
    x"60e", x"60c", x"60a", x"608", x"606", x"604", x"602", x"600", 
    x"5fd", x"5fb", x"5f9", x"5f7", x"5f5", x"5f3", x"5f1", x"5ef", 
    x"5ed", x"5eb", x"5e9", x"5e6", x"5e4", x"5e2", x"5e0", x"5de", 
    x"5dc", x"5da", x"5d7", x"5d5", x"5d3", x"5d1", x"5cf", x"5cd", 
    x"5cb", x"5c8", x"5c6", x"5c4", x"5c2", x"5c0", x"5bd", x"5bb", 
    x"5b9", x"5b7", x"5b5", x"5b3", x"5b0", x"5ae", x"5ac", x"5aa", 
    x"5a7", x"5a5", x"5a3", x"5a1", x"59f", x"59c", x"59a", x"598", 
    x"596", x"593", x"591", x"58f", x"58d", x"58a", x"588", x"586", 
    x"583", x"581", x"57f", x"57d", x"57a", x"578", x"576", x"573", 
    x"571", x"56f", x"56d", x"56a", x"568", x"566", x"563", x"561", 
    x"55f", x"55c", x"55a", x"558", x"555", x"553", x"551", x"54e", 
    x"54c", x"54a", x"547", x"545", x"543", x"540", x"53e", x"53b", 
    x"539", x"537", x"534", x"532", x"530", x"52d", x"52b", x"528", 
    x"526", x"524", x"521", x"51f", x"51c", x"51a", x"517", x"515", 
    x"513", x"510", x"50e", x"50b", x"509", x"506", x"504", x"502", 
    x"4ff", x"4fd", x"4fa", x"4f8", x"4f5", x"4f3", x"4f0", x"4ee", 
    x"4eb", x"4e9", x"4e6", x"4e4", x"4e1", x"4df", x"4dc", x"4da", 
    x"4d7", x"4d5", x"4d2", x"4d0", x"4cd", x"4cb", x"4c8", x"4c6", 
    x"4c3", x"4c1", x"4be", x"4bc", x"4b9", x"4b7", x"4b4", x"4b2", 
    x"4af", x"4ad", x"4aa", x"4a7", x"4a5", x"4a2", x"4a0", x"49d", 
    x"49b", x"498", x"496", x"493", x"490", x"48e", x"48b", x"489", 
    x"486", x"483", x"481", x"47e", x"47c", x"479", x"476", x"474", 
    x"471", x"46f", x"46c", x"469", x"467", x"464", x"462", x"45f", 
    x"45c", x"45a", x"457", x"454", x"452", x"44f", x"44c", x"44a", 
    x"447", x"444", x"442", x"43f", x"43d", x"43a", x"437", x"435", 
    x"432", x"42f", x"42c", x"42a", x"427", x"424", x"422", x"41f", 
    x"41c", x"41a", x"417", x"414", x"412", x"40f", x"40c", x"409", 
    x"407", x"404", x"401", x"3ff", x"3fc", x"3f9", x"3f6", x"3f4", 
    x"3f1", x"3ee", x"3eb", x"3e9", x"3e6", x"3e3", x"3e1", x"3de", 
    x"3db", x"3d8", x"3d6", x"3d3", x"3d0", x"3cd", x"3ca", x"3c8", 
    x"3c5", x"3c2", x"3bf", x"3bd", x"3ba", x"3b7", x"3b4", x"3b2", 
    x"3af", x"3ac", x"3a9", x"3a6", x"3a4", x"3a1", x"39e", x"39b", 
    x"398", x"396", x"393", x"390", x"38d", x"38a", x"387", x"385", 
    x"382", x"37f", x"37c", x"379", x"377", x"374", x"371", x"36e", 
    x"36b", x"368", x"366", x"363", x"360", x"35d", x"35a", x"357", 
    x"354", x"352", x"34f", x"34c", x"349", x"346", x"343", x"340", 
    x"33e", x"33b", x"338", x"335", x"332", x"32f", x"32c", x"329", 
    x"327", x"324", x"321", x"31e", x"31b", x"318", x"315", x"312", 
    x"30f", x"30c", x"30a", x"307", x"304", x"301", x"2fe", x"2fb", 
    x"2f8", x"2f5", x"2f2", x"2ef", x"2ec", x"2e9", x"2e7", x"2e4", 
    x"2e1", x"2de", x"2db", x"2d8", x"2d5", x"2d2", x"2cf", x"2cc", 
    x"2c9", x"2c6", x"2c3", x"2c0", x"2bd", x"2ba", x"2b8", x"2b5", 
    x"2b2", x"2af", x"2ac", x"2a9", x"2a6", x"2a3", x"2a0", x"29d", 
    x"29a", x"297", x"294", x"291", x"28e", x"28b", x"288", x"285", 
    x"282", x"27f", x"27c", x"279", x"276", x"273", x"270", x"26d", 
    x"26a", x"267", x"264", x"261", x"25e", x"25b", x"258", x"255", 
    x"252", x"24f", x"24c", x"249", x"246", x"243", x"240", x"23d", 
    x"23a", x"237", x"234", x"231", x"22e", x"22b", x"228", x"225", 
    x"222", x"21f", x"21c", x"219", x"216", x"213", x"210", x"20d", 
    x"20a", x"207", x"204", x"201", x"1fe", x"1fb", x"1f7", x"1f4", 
    x"1f1", x"1ee", x"1eb", x"1e8", x"1e5", x"1e2", x"1df", x"1dc", 
    x"1d9", x"1d6", x"1d3", x"1d0", x"1cd", x"1ca", x"1c7", x"1c4", 
    x"1c1", x"1bd", x"1ba", x"1b7", x"1b4", x"1b1", x"1ae", x"1ab", 
    x"1a8", x"1a5", x"1a2", x"19f", x"19c", x"199", x"196", x"192", 
    x"18f", x"18c", x"189", x"186", x"183", x"180", x"17d", x"17a", 
    x"177", x"174", x"171", x"16d", x"16a", x"167", x"164", x"161", 
    x"15e", x"15b", x"158", x"155", x"152", x"14e", x"14b", x"148", 
    x"145", x"142", x"13f", x"13c", x"139", x"136", x"133", x"12f", 
    x"12c", x"129", x"126", x"123", x"120", x"11d", x"11a", x"117", 
    x"113", x"110", x"10d", x"10a", x"107", x"104", x"101", x"0fe", 
    x"0fb", x"0f7", x"0f4", x"0f1", x"0ee", x"0eb", x"0e8", x"0e5", 
    x"0e2", x"0df", x"0db", x"0d8", x"0d5", x"0d2", x"0cf", x"0cc", 
    x"0c9", x"0c6", x"0c2", x"0bf", x"0bc", x"0b9", x"0b6", x"0b3", 
    x"0b0", x"0ac", x"0a9", x"0a6", x"0a3", x"0a0", x"09d", x"09a", 
    x"097", x"093", x"090", x"08d", x"08a", x"087", x"084", x"081", 
    x"07e", x"07a", x"077", x"074", x"071", x"06e", x"06b", x"068", 
    x"064", x"061", x"05e", x"05b", x"058", x"055", x"052", x"04e", 
    x"04b", x"048", x"045", x"042", x"03f", x"03c", x"039", x"035", 
    x"032", x"02f", x"02c", x"029", x"026", x"023", x"01f", x"01c", 
    x"019", x"016", x"013", x"010", x"00d", x"009", x"006", x"003", 
    x"000", x"ffd", x"ffa", x"ff7", x"ff3", x"ff0", x"fed", x"fea", 
    x"fe7", x"fe4", x"fe1", x"fdd", x"fda", x"fd7", x"fd4", x"fd1", 
    x"fce", x"fcb", x"fc7", x"fc4", x"fc1", x"fbe", x"fbb", x"fb8", 
    x"fb5", x"fb2", x"fae", x"fab", x"fa8", x"fa5", x"fa2", x"f9f", 
    x"f9c", x"f98", x"f95", x"f92", x"f8f", x"f8c", x"f89", x"f86", 
    x"f82", x"f7f", x"f7c", x"f79", x"f76", x"f73", x"f70", x"f6d", 
    x"f69", x"f66", x"f63", x"f60", x"f5d", x"f5a", x"f57", x"f54", 
    x"f50", x"f4d", x"f4a", x"f47", x"f44", x"f41", x"f3e", x"f3a", 
    x"f37", x"f34", x"f31", x"f2e", x"f2b", x"f28", x"f25", x"f21", 
    x"f1e", x"f1b", x"f18", x"f15", x"f12", x"f0f", x"f0c", x"f09", 
    x"f05", x"f02", x"eff", x"efc", x"ef9", x"ef6", x"ef3", x"ef0", 
    x"eed", x"ee9", x"ee6", x"ee3", x"ee0", x"edd", x"eda", x"ed7", 
    x"ed4", x"ed1", x"ecd", x"eca", x"ec7", x"ec4", x"ec1", x"ebe", 
    x"ebb", x"eb8", x"eb5", x"eb2", x"eae", x"eab", x"ea8", x"ea5", 
    x"ea2", x"e9f", x"e9c", x"e99", x"e96", x"e93", x"e8f", x"e8c", 
    x"e89", x"e86", x"e83", x"e80", x"e7d", x"e7a", x"e77", x"e74", 
    x"e71", x"e6e", x"e6a", x"e67", x"e64", x"e61", x"e5e", x"e5b", 
    x"e58", x"e55", x"e52", x"e4f", x"e4c", x"e49", x"e46", x"e43", 
    x"e3f", x"e3c", x"e39", x"e36", x"e33", x"e30", x"e2d", x"e2a", 
    x"e27", x"e24", x"e21", x"e1e", x"e1b", x"e18", x"e15", x"e12", 
    x"e0f", x"e0c", x"e09", x"e05", x"e02", x"dff", x"dfc", x"df9", 
    x"df6", x"df3", x"df0", x"ded", x"dea", x"de7", x"de4", x"de1", 
    x"dde", x"ddb", x"dd8", x"dd5", x"dd2", x"dcf", x"dcc", x"dc9", 
    x"dc6", x"dc3", x"dc0", x"dbd", x"dba", x"db7", x"db4", x"db1", 
    x"dae", x"dab", x"da8", x"da5", x"da2", x"d9f", x"d9c", x"d99", 
    x"d96", x"d93", x"d90", x"d8d", x"d8a", x"d87", x"d84", x"d81", 
    x"d7e", x"d7b", x"d78", x"d75", x"d72", x"d6f", x"d6c", x"d69", 
    x"d66", x"d63", x"d60", x"d5d", x"d5a", x"d57", x"d54", x"d51", 
    x"d4e", x"d4b", x"d48", x"d46", x"d43", x"d40", x"d3d", x"d3a", 
    x"d37", x"d34", x"d31", x"d2e", x"d2b", x"d28", x"d25", x"d22", 
    x"d1f", x"d1c", x"d19", x"d17", x"d14", x"d11", x"d0e", x"d0b", 
    x"d08", x"d05", x"d02", x"cff", x"cfc", x"cf9", x"cf6", x"cf4", 
    x"cf1", x"cee", x"ceb", x"ce8", x"ce5", x"ce2", x"cdf", x"cdc", 
    x"cd9", x"cd7", x"cd4", x"cd1", x"cce", x"ccb", x"cc8", x"cc5", 
    x"cc2", x"cc0", x"cbd", x"cba", x"cb7", x"cb4", x"cb1", x"cae", 
    x"cac", x"ca9", x"ca6", x"ca3", x"ca0", x"c9d", x"c9a", x"c98", 
    x"c95", x"c92", x"c8f", x"c8c", x"c89", x"c87", x"c84", x"c81", 
    x"c7e", x"c7b", x"c79", x"c76", x"c73", x"c70", x"c6d", x"c6a", 
    x"c68", x"c65", x"c62", x"c5f", x"c5c", x"c5a", x"c57", x"c54", 
    x"c51", x"c4e", x"c4c", x"c49", x"c46", x"c43", x"c41", x"c3e", 
    x"c3b", x"c38", x"c36", x"c33", x"c30", x"c2d", x"c2a", x"c28", 
    x"c25", x"c22", x"c1f", x"c1d", x"c1a", x"c17", x"c15", x"c12", 
    x"c0f", x"c0c", x"c0a", x"c07", x"c04", x"c01", x"bff", x"bfc", 
    x"bf9", x"bf7", x"bf4", x"bf1", x"bee", x"bec", x"be9", x"be6", 
    x"be4", x"be1", x"bde", x"bdc", x"bd9", x"bd6", x"bd4", x"bd1", 
    x"bce", x"bcb", x"bc9", x"bc6", x"bc3", x"bc1", x"bbe", x"bbc", 
    x"bb9", x"bb6", x"bb4", x"bb1", x"bae", x"bac", x"ba9", x"ba6", 
    x"ba4", x"ba1", x"b9e", x"b9c", x"b99", x"b97", x"b94", x"b91", 
    x"b8f", x"b8c", x"b8a", x"b87", x"b84", x"b82", x"b7f", x"b7d", 
    x"b7a", x"b77", x"b75", x"b72", x"b70", x"b6d", x"b6a", x"b68", 
    x"b65", x"b63", x"b60", x"b5e", x"b5b", x"b59", x"b56", x"b53", 
    x"b51", x"b4e", x"b4c", x"b49", x"b47", x"b44", x"b42", x"b3f", 
    x"b3d", x"b3a", x"b38", x"b35", x"b33", x"b30", x"b2e", x"b2b", 
    x"b29", x"b26", x"b24", x"b21", x"b1f", x"b1c", x"b1a", x"b17", 
    x"b15", x"b12", x"b10", x"b0d", x"b0b", x"b08", x"b06", x"b03", 
    x"b01", x"afe", x"afc", x"afa", x"af7", x"af5", x"af2", x"af0", 
    x"aed", x"aeb", x"ae9", x"ae6", x"ae4", x"ae1", x"adf", x"adc", 
    x"ada", x"ad8", x"ad5", x"ad3", x"ad0", x"ace", x"acc", x"ac9", 
    x"ac7", x"ac5", x"ac2", x"ac0", x"abd", x"abb", x"ab9", x"ab6", 
    x"ab4", x"ab2", x"aaf", x"aad", x"aab", x"aa8", x"aa6", x"aa4", 
    x"aa1", x"a9f", x"a9d", x"a9a", x"a98", x"a96", x"a93", x"a91", 
    x"a8f", x"a8d", x"a8a", x"a88", x"a86", x"a83", x"a81", x"a7f", 
    x"a7d", x"a7a", x"a78", x"a76", x"a73", x"a71", x"a6f", x"a6d", 
    x"a6a", x"a68", x"a66", x"a64", x"a61", x"a5f", x"a5d", x"a5b", 
    x"a59", x"a56", x"a54", x"a52", x"a50", x"a4d", x"a4b", x"a49", 
    x"a47", x"a45", x"a43", x"a40", x"a3e", x"a3c", x"a3a", x"a38", 
    x"a35", x"a33", x"a31", x"a2f", x"a2d", x"a2b", x"a29", x"a26", 
    x"a24", x"a22", x"a20", x"a1e", x"a1c", x"a1a", x"a17", x"a15", 
    x"a13", x"a11", x"a0f", x"a0d", x"a0b", x"a09", x"a07", x"a05", 
    x"a03", x"a00", x"9fe", x"9fc", x"9fa", x"9f8", x"9f6", x"9f4", 
    x"9f2", x"9f0", x"9ee", x"9ec", x"9ea", x"9e8", x"9e6", x"9e4", 
    x"9e2", x"9e0", x"9de", x"9dc", x"9da", x"9d8", x"9d6", x"9d4", 
    x"9d2", x"9d0", x"9ce", x"9cc", x"9ca", x"9c8", x"9c6", x"9c4", 
    x"9c2", x"9c0", x"9be", x"9bc", x"9ba", x"9b8", x"9b6", x"9b4", 
    x"9b2", x"9b0", x"9ae", x"9ac", x"9ab", x"9a9", x"9a7", x"9a5", 
    x"9a3", x"9a1", x"99f", x"99d", x"99b", x"999", x"998", x"996", 
    x"994", x"992", x"990", x"98e", x"98c", x"98b", x"989", x"987", 
    x"985", x"983", x"981", x"97f", x"97e", x"97c", x"97a", x"978", 
    x"976", x"975", x"973", x"971", x"96f", x"96d", x"96c", x"96a", 
    x"968", x"966", x"965", x"963", x"961", x"95f", x"95d", x"95c", 
    x"95a", x"958", x"957", x"955", x"953", x"951", x"950", x"94e", 
    x"94c", x"94a", x"949", x"947", x"945", x"944", x"942", x"940", 
    x"93f", x"93d", x"93b", x"93a", x"938", x"936", x"935", x"933", 
    x"931", x"930", x"92e", x"92c", x"92b", x"929", x"927", x"926", 
    x"924", x"923", x"921", x"91f", x"91e", x"91c", x"91b", x"919", 
    x"917", x"916", x"914", x"913", x"911", x"910", x"90e", x"90c", 
    x"90b", x"909", x"908", x"906", x"905", x"903", x"902", x"900", 
    x"8ff", x"8fd", x"8fc", x"8fa", x"8f9", x"8f7", x"8f6", x"8f4", 
    x"8f3", x"8f1", x"8f0", x"8ee", x"8ed", x"8eb", x"8ea", x"8e8", 
    x"8e7", x"8e6", x"8e4", x"8e3", x"8e1", x"8e0", x"8de", x"8dd", 
    x"8dc", x"8da", x"8d9", x"8d7", x"8d6", x"8d5", x"8d3", x"8d2", 
    x"8d0", x"8cf", x"8ce", x"8cc", x"8cb", x"8ca", x"8c8", x"8c7", 
    x"8c6", x"8c4", x"8c3", x"8c2", x"8c0", x"8bf", x"8be", x"8bc", 
    x"8bb", x"8ba", x"8b8", x"8b7", x"8b6", x"8b4", x"8b3", x"8b2", 
    x"8b1", x"8af", x"8ae", x"8ad", x"8ac", x"8aa", x"8a9", x"8a8", 
    x"8a7", x"8a5", x"8a4", x"8a3", x"8a2", x"8a0", x"89f", x"89e", 
    x"89d", x"89c", x"89a", x"899", x"898", x"897", x"896", x"895", 
    x"893", x"892", x"891", x"890", x"88f", x"88e", x"88c", x"88b", 
    x"88a", x"889", x"888", x"887", x"886", x"885", x"883", x"882", 
    x"881", x"880", x"87f", x"87e", x"87d", x"87c", x"87b", x"87a", 
    x"879", x"878", x"877", x"876", x"874", x"873", x"872", x"871", 
    x"870", x"86f", x"86e", x"86d", x"86c", x"86b", x"86a", x"869", 
    x"868", x"867", x"866", x"865", x"864", x"863", x"862", x"862", 
    x"861", x"860", x"85f", x"85e", x"85d", x"85c", x"85b", x"85a", 
    x"859", x"858", x"857", x"856", x"856", x"855", x"854", x"853", 
    x"852", x"851", x"850", x"84f", x"84f", x"84e", x"84d", x"84c", 
    x"84b", x"84a", x"849", x"849", x"848", x"847", x"846", x"845", 
    x"845", x"844", x"843", x"842", x"841", x"841", x"840", x"83f", 
    x"83e", x"83e", x"83d", x"83c", x"83b", x"83b", x"83a", x"839", 
    x"838", x"838", x"837", x"836", x"836", x"835", x"834", x"833", 
    x"833", x"832", x"831", x"831", x"830", x"82f", x"82f", x"82e", 
    x"82d", x"82d", x"82c", x"82b", x"82b", x"82a", x"82a", x"829", 
    x"828", x"828", x"827", x"827", x"826", x"825", x"825", x"824", 
    x"824", x"823", x"822", x"822", x"821", x"821", x"820", x"820", 
    x"81f", x"81f", x"81e", x"81e", x"81d", x"81d", x"81c", x"81b", 
    x"81b", x"81a", x"81a", x"81a", x"819", x"819", x"818", x"818", 
    x"817", x"817", x"816", x"816", x"815", x"815", x"814", x"814", 
    x"814", x"813", x"813", x"812", x"812", x"812", x"811", x"811", 
    x"810", x"810", x"810", x"80f", x"80f", x"80f", x"80e", x"80e", 
    x"80d", x"80d", x"80d", x"80c", x"80c", x"80c", x"80b", x"80b", 
    x"80b", x"80b", x"80a", x"80a", x"80a", x"809", x"809", x"809", 
    x"809", x"808", x"808", x"808", x"808", x"807", x"807", x"807", 
    x"807", x"806", x"806", x"806", x"806", x"805", x"805", x"805", 
    x"805", x"805", x"804", x"804", x"804", x"804", x"804", x"804", 
    x"803", x"803", x"803", x"803", x"803", x"803", x"803", x"803", 
    x"802", x"802", x"802", x"802", x"802", x"802", x"802", x"802", 
    x"802", x"802", x"801", x"801", x"801", x"801", x"801", x"801", 
    x"801", x"801", x"801", x"801", x"801", x"801", x"801", x"801", 
    x"801", x"801", x"801", x"801", x"801", x"801", x"801", x"801", 
    x"801", x"801", x"801", x"801", x"801", x"801", x"801", x"802", 
    x"802", x"802", x"802", x"802", x"802", x"802", x"802", x"802", 
    x"802", x"803", x"803", x"803", x"803", x"803", x"803", x"803", 
    x"803", x"804", x"804", x"804", x"804", x"804", x"804", x"805", 
    x"805", x"805", x"805", x"805", x"806", x"806", x"806", x"806", 
    x"807", x"807", x"807", x"807", x"808", x"808", x"808", x"808", 
    x"809", x"809", x"809", x"809", x"80a", x"80a", x"80a", x"80b", 
    x"80b", x"80b", x"80b", x"80c", x"80c", x"80c", x"80d", x"80d", 
    x"80d", x"80e", x"80e", x"80f", x"80f", x"80f", x"810", x"810", 
    x"810", x"811", x"811", x"812", x"812", x"812", x"813", x"813", 
    x"814", x"814", x"814", x"815", x"815", x"816", x"816", x"817", 
    x"817", x"818", x"818", x"819", x"819", x"81a", x"81a", x"81a", 
    x"81b", x"81b", x"81c", x"81d", x"81d", x"81e", x"81e", x"81f", 
    x"81f", x"820", x"820", x"821", x"821", x"822", x"822", x"823", 
    x"824", x"824", x"825", x"825", x"826", x"827", x"827", x"828", 
    x"828", x"829", x"82a", x"82a", x"82b", x"82b", x"82c", x"82d", 
    x"82d", x"82e", x"82f", x"82f", x"830", x"831", x"831", x"832", 
    x"833", x"833", x"834", x"835", x"836", x"836", x"837", x"838", 
    x"838", x"839", x"83a", x"83b", x"83b", x"83c", x"83d", x"83e", 
    x"83e", x"83f", x"840", x"841", x"841", x"842", x"843", x"844", 
    x"845", x"845", x"846", x"847", x"848", x"849", x"849", x"84a", 
    x"84b", x"84c", x"84d", x"84e", x"84f", x"84f", x"850", x"851", 
    x"852", x"853", x"854", x"855", x"856", x"856", x"857", x"858", 
    x"859", x"85a", x"85b", x"85c", x"85d", x"85e", x"85f", x"860", 
    x"861", x"862", x"862", x"863", x"864", x"865", x"866", x"867", 
    x"868", x"869", x"86a", x"86b", x"86c", x"86d", x"86e", x"86f", 
    x"870", x"871", x"872", x"873", x"874", x"876", x"877", x"878", 
    x"879", x"87a", x"87b", x"87c", x"87d", x"87e", x"87f", x"880", 
    x"881", x"882", x"883", x"885", x"886", x"887", x"888", x"889", 
    x"88a", x"88b", x"88c", x"88e", x"88f", x"890", x"891", x"892", 
    x"893", x"895", x"896", x"897", x"898", x"899", x"89a", x"89c", 
    x"89d", x"89e", x"89f", x"8a0", x"8a2", x"8a3", x"8a4", x"8a5", 
    x"8a7", x"8a8", x"8a9", x"8aa", x"8ac", x"8ad", x"8ae", x"8af", 
    x"8b1", x"8b2", x"8b3", x"8b4", x"8b6", x"8b7", x"8b8", x"8ba", 
    x"8bb", x"8bc", x"8be", x"8bf", x"8c0", x"8c2", x"8c3", x"8c4", 
    x"8c6", x"8c7", x"8c8", x"8ca", x"8cb", x"8cc", x"8ce", x"8cf", 
    x"8d0", x"8d2", x"8d3", x"8d5", x"8d6", x"8d7", x"8d9", x"8da", 
    x"8dc", x"8dd", x"8de", x"8e0", x"8e1", x"8e3", x"8e4", x"8e6", 
    x"8e7", x"8e8", x"8ea", x"8eb", x"8ed", x"8ee", x"8f0", x"8f1", 
    x"8f3", x"8f4", x"8f6", x"8f7", x"8f9", x"8fa", x"8fc", x"8fd", 
    x"8ff", x"900", x"902", x"903", x"905", x"906", x"908", x"909", 
    x"90b", x"90c", x"90e", x"910", x"911", x"913", x"914", x"916", 
    x"917", x"919", x"91b", x"91c", x"91e", x"91f", x"921", x"923", 
    x"924", x"926", x"927", x"929", x"92b", x"92c", x"92e", x"930", 
    x"931", x"933", x"935", x"936", x"938", x"93a", x"93b", x"93d", 
    x"93f", x"940", x"942", x"944", x"945", x"947", x"949", x"94a", 
    x"94c", x"94e", x"950", x"951", x"953", x"955", x"957", x"958", 
    x"95a", x"95c", x"95d", x"95f", x"961", x"963", x"965", x"966", 
    x"968", x"96a", x"96c", x"96d", x"96f", x"971", x"973", x"975", 
    x"976", x"978", x"97a", x"97c", x"97e", x"97f", x"981", x"983", 
    x"985", x"987", x"989", x"98b", x"98c", x"98e", x"990", x"992", 
    x"994", x"996", x"998", x"999", x"99b", x"99d", x"99f", x"9a1", 
    x"9a3", x"9a5", x"9a7", x"9a9", x"9ab", x"9ac", x"9ae", x"9b0", 
    x"9b2", x"9b4", x"9b6", x"9b8", x"9ba", x"9bc", x"9be", x"9c0", 
    x"9c2", x"9c4", x"9c6", x"9c8", x"9ca", x"9cc", x"9ce", x"9d0", 
    x"9d2", x"9d4", x"9d6", x"9d8", x"9da", x"9dc", x"9de", x"9e0", 
    x"9e2", x"9e4", x"9e6", x"9e8", x"9ea", x"9ec", x"9ee", x"9f0", 
    x"9f2", x"9f4", x"9f6", x"9f8", x"9fa", x"9fc", x"9fe", x"a00", 
    x"a03", x"a05", x"a07", x"a09", x"a0b", x"a0d", x"a0f", x"a11", 
    x"a13", x"a15", x"a17", x"a1a", x"a1c", x"a1e", x"a20", x"a22", 
    x"a24", x"a26", x"a29", x"a2b", x"a2d", x"a2f", x"a31", x"a33", 
    x"a35", x"a38", x"a3a", x"a3c", x"a3e", x"a40", x"a43", x"a45", 
    x"a47", x"a49", x"a4b", x"a4d", x"a50", x"a52", x"a54", x"a56", 
    x"a59", x"a5b", x"a5d", x"a5f", x"a61", x"a64", x"a66", x"a68", 
    x"a6a", x"a6d", x"a6f", x"a71", x"a73", x"a76", x"a78", x"a7a", 
    x"a7d", x"a7f", x"a81", x"a83", x"a86", x"a88", x"a8a", x"a8d", 
    x"a8f", x"a91", x"a93", x"a96", x"a98", x"a9a", x"a9d", x"a9f", 
    x"aa1", x"aa4", x"aa6", x"aa8", x"aab", x"aad", x"aaf", x"ab2", 
    x"ab4", x"ab6", x"ab9", x"abb", x"abd", x"ac0", x"ac2", x"ac5", 
    x"ac7", x"ac9", x"acc", x"ace", x"ad0", x"ad3", x"ad5", x"ad8", 
    x"ada", x"adc", x"adf", x"ae1", x"ae4", x"ae6", x"ae9", x"aeb", 
    x"aed", x"af0", x"af2", x"af5", x"af7", x"afa", x"afc", x"afe", 
    x"b01", x"b03", x"b06", x"b08", x"b0b", x"b0d", x"b10", x"b12", 
    x"b15", x"b17", x"b1a", x"b1c", x"b1f", x"b21", x"b24", x"b26", 
    x"b29", x"b2b", x"b2e", x"b30", x"b33", x"b35", x"b38", x"b3a", 
    x"b3d", x"b3f", x"b42", x"b44", x"b47", x"b49", x"b4c", x"b4e", 
    x"b51", x"b53", x"b56", x"b59", x"b5b", x"b5e", x"b60", x"b63", 
    x"b65", x"b68", x"b6a", x"b6d", x"b70", x"b72", x"b75", x"b77", 
    x"b7a", x"b7d", x"b7f", x"b82", x"b84", x"b87", x"b8a", x"b8c", 
    x"b8f", x"b91", x"b94", x"b97", x"b99", x"b9c", x"b9e", x"ba1", 
    x"ba4", x"ba6", x"ba9", x"bac", x"bae", x"bb1", x"bb4", x"bb6", 
    x"bb9", x"bbc", x"bbe", x"bc1", x"bc3", x"bc6", x"bc9", x"bcb", 
    x"bce", x"bd1", x"bd4", x"bd6", x"bd9", x"bdc", x"bde", x"be1", 
    x"be4", x"be6", x"be9", x"bec", x"bee", x"bf1", x"bf4", x"bf7", 
    x"bf9", x"bfc", x"bff", x"c01", x"c04", x"c07", x"c0a", x"c0c", 
    x"c0f", x"c12", x"c15", x"c17", x"c1a", x"c1d", x"c1f", x"c22", 
    x"c25", x"c28", x"c2a", x"c2d", x"c30", x"c33", x"c36", x"c38", 
    x"c3b", x"c3e", x"c41", x"c43", x"c46", x"c49", x"c4c", x"c4e", 
    x"c51", x"c54", x"c57", x"c5a", x"c5c", x"c5f", x"c62", x"c65", 
    x"c68", x"c6a", x"c6d", x"c70", x"c73", x"c76", x"c79", x"c7b", 
    x"c7e", x"c81", x"c84", x"c87", x"c89", x"c8c", x"c8f", x"c92", 
    x"c95", x"c98", x"c9a", x"c9d", x"ca0", x"ca3", x"ca6", x"ca9", 
    x"cac", x"cae", x"cb1", x"cb4", x"cb7", x"cba", x"cbd", x"cc0", 
    x"cc2", x"cc5", x"cc8", x"ccb", x"cce", x"cd1", x"cd4", x"cd7", 
    x"cd9", x"cdc", x"cdf", x"ce2", x"ce5", x"ce8", x"ceb", x"cee", 
    x"cf1", x"cf4", x"cf6", x"cf9", x"cfc", x"cff", x"d02", x"d05", 
    x"d08", x"d0b", x"d0e", x"d11", x"d14", x"d17", x"d19", x"d1c", 
    x"d1f", x"d22", x"d25", x"d28", x"d2b", x"d2e", x"d31", x"d34", 
    x"d37", x"d3a", x"d3d", x"d40", x"d43", x"d46", x"d48", x"d4b", 
    x"d4e", x"d51", x"d54", x"d57", x"d5a", x"d5d", x"d60", x"d63", 
    x"d66", x"d69", x"d6c", x"d6f", x"d72", x"d75", x"d78", x"d7b", 
    x"d7e", x"d81", x"d84", x"d87", x"d8a", x"d8d", x"d90", x"d93", 
    x"d96", x"d99", x"d9c", x"d9f", x"da2", x"da5", x"da8", x"dab", 
    x"dae", x"db1", x"db4", x"db7", x"dba", x"dbd", x"dc0", x"dc3", 
    x"dc6", x"dc9", x"dcc", x"dcf", x"dd2", x"dd5", x"dd8", x"ddb", 
    x"dde", x"de1", x"de4", x"de7", x"dea", x"ded", x"df0", x"df3", 
    x"df6", x"df9", x"dfc", x"dff", x"e02", x"e05", x"e09", x"e0c", 
    x"e0f", x"e12", x"e15", x"e18", x"e1b", x"e1e", x"e21", x"e24", 
    x"e27", x"e2a", x"e2d", x"e30", x"e33", x"e36", x"e39", x"e3c", 
    x"e3f", x"e43", x"e46", x"e49", x"e4c", x"e4f", x"e52", x"e55", 
    x"e58", x"e5b", x"e5e", x"e61", x"e64", x"e67", x"e6a", x"e6e", 
    x"e71", x"e74", x"e77", x"e7a", x"e7d", x"e80", x"e83", x"e86", 
    x"e89", x"e8c", x"e8f", x"e93", x"e96", x"e99", x"e9c", x"e9f", 
    x"ea2", x"ea5", x"ea8", x"eab", x"eae", x"eb2", x"eb5", x"eb8", 
    x"ebb", x"ebe", x"ec1", x"ec4", x"ec7", x"eca", x"ecd", x"ed1", 
    x"ed4", x"ed7", x"eda", x"edd", x"ee0", x"ee3", x"ee6", x"ee9", 
    x"eed", x"ef0", x"ef3", x"ef6", x"ef9", x"efc", x"eff", x"f02", 
    x"f05", x"f09", x"f0c", x"f0f", x"f12", x"f15", x"f18", x"f1b", 
    x"f1e", x"f21", x"f25", x"f28", x"f2b", x"f2e", x"f31", x"f34", 
    x"f37", x"f3a", x"f3e", x"f41", x"f44", x"f47", x"f4a", x"f4d", 
    x"f50", x"f54", x"f57", x"f5a", x"f5d", x"f60", x"f63", x"f66", 
    x"f69", x"f6d", x"f70", x"f73", x"f76", x"f79", x"f7c", x"f7f", 
    x"f82", x"f86", x"f89", x"f8c", x"f8f", x"f92", x"f95", x"f98", 
    x"f9c", x"f9f", x"fa2", x"fa5", x"fa8", x"fab", x"fae", x"fb2", 
    x"fb5", x"fb8", x"fbb", x"fbe", x"fc1", x"fc4", x"fc7", x"fcb", 
    x"fce", x"fd1", x"fd4", x"fd7", x"fda", x"fdd", x"fe1", x"fe4", 
    x"fe7", x"fea", x"fed", x"ff0", x"ff3", x"ff7", x"ffa", x"ffd", 
    x"000", x"003", x"006", x"009", x"00d", x"010", x"013", x"016", 
    x"019", x"01c", x"01f", x"023", x"026", x"029", x"02c", x"02f", 
    x"032", x"035", x"039", x"03c", x"03f", x"042", x"045", x"048", 
    x"04b", x"04e", x"052", x"055", x"058", x"05b", x"05e", x"061", 
    x"064", x"068", x"06b", x"06e", x"071", x"074", x"077", x"07a", 
    x"07e", x"081", x"084", x"087", x"08a", x"08d", x"090", x"093", 
    x"097", x"09a", x"09d", x"0a0", x"0a3", x"0a6", x"0a9", x"0ac", 
    x"0b0", x"0b3", x"0b6", x"0b9", x"0bc", x"0bf", x"0c2", x"0c6", 
    x"0c9", x"0cc", x"0cf", x"0d2", x"0d5", x"0d8", x"0db", x"0df", 
    x"0e2", x"0e5", x"0e8", x"0eb", x"0ee", x"0f1", x"0f4", x"0f7", 
    x"0fb", x"0fe", x"101", x"104", x"107", x"10a", x"10d", x"110", 
    x"113", x"117", x"11a", x"11d", x"120", x"123", x"126", x"129", 
    x"12c", x"12f", x"133", x"136", x"139", x"13c", x"13f", x"142", 
    x"145", x"148", x"14b", x"14e", x"152", x"155", x"158", x"15b", 
    x"15e", x"161", x"164", x"167", x"16a", x"16d", x"171", x"174", 
    x"177", x"17a", x"17d", x"180", x"183", x"186", x"189", x"18c", 
    x"18f", x"192", x"196", x"199", x"19c", x"19f", x"1a2", x"1a5", 
    x"1a8", x"1ab", x"1ae", x"1b1", x"1b4", x"1b7", x"1ba", x"1bd", 
    x"1c1", x"1c4", x"1c7", x"1ca", x"1cd", x"1d0", x"1d3", x"1d6", 
    x"1d9", x"1dc", x"1df", x"1e2", x"1e5", x"1e8", x"1eb", x"1ee", 
    x"1f1", x"1f4", x"1f7", x"1fb", x"1fe", x"201", x"204", x"207", 
    x"20a", x"20d", x"210", x"213", x"216", x"219", x"21c", x"21f", 
    x"222", x"225", x"228", x"22b", x"22e", x"231", x"234", x"237", 
    x"23a", x"23d", x"240", x"243", x"246", x"249", x"24c", x"24f", 
    x"252", x"255", x"258", x"25b", x"25e", x"261", x"264", x"267", 
    x"26a", x"26d", x"270", x"273", x"276", x"279", x"27c", x"27f", 
    x"282", x"285", x"288", x"28b", x"28e", x"291", x"294", x"297", 
    x"29a", x"29d", x"2a0", x"2a3", x"2a6", x"2a9", x"2ac", x"2af", 
    x"2b2", x"2b5", x"2b8", x"2ba", x"2bd", x"2c0", x"2c3", x"2c6", 
    x"2c9", x"2cc", x"2cf", x"2d2", x"2d5", x"2d8", x"2db", x"2de", 
    x"2e1", x"2e4", x"2e7", x"2e9", x"2ec", x"2ef", x"2f2", x"2f5", 
    x"2f8", x"2fb", x"2fe", x"301", x"304", x"307", x"30a", x"30c", 
    x"30f", x"312", x"315", x"318", x"31b", x"31e", x"321", x"324", 
    x"327", x"329", x"32c", x"32f", x"332", x"335", x"338", x"33b", 
    x"33e", x"340", x"343", x"346", x"349", x"34c", x"34f", x"352", 
    x"354", x"357", x"35a", x"35d", x"360", x"363", x"366", x"368", 
    x"36b", x"36e", x"371", x"374", x"377", x"379", x"37c", x"37f", 
    x"382", x"385", x"387", x"38a", x"38d", x"390", x"393", x"396", 
    x"398", x"39b", x"39e", x"3a1", x"3a4", x"3a6", x"3a9", x"3ac", 
    x"3af", x"3b2", x"3b4", x"3b7", x"3ba", x"3bd", x"3bf", x"3c2", 
    x"3c5", x"3c8", x"3ca", x"3cd", x"3d0", x"3d3", x"3d6", x"3d8", 
    x"3db", x"3de", x"3e1", x"3e3", x"3e6", x"3e9", x"3eb", x"3ee", 
    x"3f1", x"3f4", x"3f6", x"3f9", x"3fc", x"3ff", x"401", x"404", 
    x"407", x"409", x"40c", x"40f", x"412", x"414", x"417", x"41a", 
    x"41c", x"41f", x"422", x"424", x"427", x"42a", x"42c", x"42f", 
    x"432", x"435", x"437", x"43a", x"43d", x"43f", x"442", x"444", 
    x"447", x"44a", x"44c", x"44f", x"452", x"454", x"457", x"45a", 
    x"45c", x"45f", x"462", x"464", x"467", x"469", x"46c", x"46f", 
    x"471", x"474", x"476", x"479", x"47c", x"47e", x"481", x"483", 
    x"486", x"489", x"48b", x"48e", x"490", x"493", x"496", x"498", 
    x"49b", x"49d", x"4a0", x"4a2", x"4a5", x"4a7", x"4aa", x"4ad", 
    x"4af", x"4b2", x"4b4", x"4b7", x"4b9", x"4bc", x"4be", x"4c1", 
    x"4c3", x"4c6", x"4c8", x"4cb", x"4cd", x"4d0", x"4d2", x"4d5", 
    x"4d7", x"4da", x"4dc", x"4df", x"4e1", x"4e4", x"4e6", x"4e9", 
    x"4eb", x"4ee", x"4f0", x"4f3", x"4f5", x"4f8", x"4fa", x"4fd", 
    x"4ff", x"502", x"504", x"506", x"509", x"50b", x"50e", x"510", 
    x"513", x"515", x"517", x"51a", x"51c", x"51f", x"521", x"524", 
    x"526", x"528", x"52b", x"52d", x"530", x"532", x"534", x"537", 
    x"539", x"53b", x"53e", x"540", x"543", x"545", x"547", x"54a", 
    x"54c", x"54e", x"551", x"553", x"555", x"558", x"55a", x"55c", 
    x"55f", x"561", x"563", x"566", x"568", x"56a", x"56d", x"56f", 
    x"571", x"573", x"576", x"578", x"57a", x"57d", x"57f", x"581", 
    x"583", x"586", x"588", x"58a", x"58d", x"58f", x"591", x"593", 
    x"596", x"598", x"59a", x"59c", x"59f", x"5a1", x"5a3", x"5a5", 
    x"5a7", x"5aa", x"5ac", x"5ae", x"5b0", x"5b3", x"5b5", x"5b7", 
    x"5b9", x"5bb", x"5bd", x"5c0", x"5c2", x"5c4", x"5c6", x"5c8", 
    x"5cb", x"5cd", x"5cf", x"5d1", x"5d3", x"5d5", x"5d7", x"5da", 
    x"5dc", x"5de", x"5e0", x"5e2", x"5e4", x"5e6", x"5e9", x"5eb", 
    x"5ed", x"5ef", x"5f1", x"5f3", x"5f5", x"5f7", x"5f9", x"5fb", 
    x"5fd", x"600", x"602", x"604", x"606", x"608", x"60a", x"60c", 
    x"60e", x"610", x"612", x"614", x"616", x"618", x"61a", x"61c", 
    x"61e", x"620", x"622", x"624", x"626", x"628", x"62a", x"62c", 
    x"62e", x"630", x"632", x"634", x"636", x"638", x"63a", x"63c", 
    x"63e", x"640", x"642", x"644", x"646", x"648", x"64a", x"64c", 
    x"64e", x"650", x"652", x"654", x"655", x"657", x"659", x"65b", 
    x"65d", x"65f", x"661", x"663", x"665", x"667", x"668", x"66a", 
    x"66c", x"66e", x"670", x"672", x"674", x"675", x"677", x"679", 
    x"67b", x"67d", x"67f", x"681", x"682", x"684", x"686", x"688", 
    x"68a", x"68b", x"68d", x"68f", x"691", x"693", x"694", x"696", 
    x"698", x"69a", x"69b", x"69d", x"69f", x"6a1", x"6a3", x"6a4", 
    x"6a6", x"6a8", x"6a9", x"6ab", x"6ad", x"6af", x"6b0", x"6b2", 
    x"6b4", x"6b6", x"6b7", x"6b9", x"6bb", x"6bc", x"6be", x"6c0", 
    x"6c1", x"6c3", x"6c5", x"6c6", x"6c8", x"6ca", x"6cb", x"6cd", 
    x"6cf", x"6d0", x"6d2", x"6d4", x"6d5", x"6d7", x"6d9", x"6da", 
    x"6dc", x"6dd", x"6df", x"6e1", x"6e2", x"6e4", x"6e5", x"6e7", 
    x"6e9", x"6ea", x"6ec", x"6ed", x"6ef", x"6f0", x"6f2", x"6f4", 
    x"6f5", x"6f7", x"6f8", x"6fa", x"6fb", x"6fd", x"6fe", x"700", 
    x"701", x"703", x"704", x"706", x"707", x"709", x"70a", x"70c", 
    x"70d", x"70f", x"710", x"712", x"713", x"715", x"716", x"718", 
    x"719", x"71a", x"71c", x"71d", x"71f", x"720", x"722", x"723", 
    x"724", x"726", x"727", x"729", x"72a", x"72b", x"72d", x"72e", 
    x"730", x"731", x"732", x"734", x"735", x"736", x"738", x"739", 
    x"73a", x"73c", x"73d", x"73e", x"740", x"741", x"742", x"744", 
    x"745", x"746", x"748", x"749", x"74a", x"74c", x"74d", x"74e", 
    x"74f", x"751", x"752", x"753", x"754", x"756", x"757", x"758", 
    x"759", x"75b", x"75c", x"75d", x"75e", x"760", x"761", x"762", 
    x"763", x"764", x"766", x"767", x"768", x"769", x"76a", x"76b", 
    x"76d", x"76e", x"76f", x"770", x"771", x"772", x"774", x"775", 
    x"776", x"777", x"778", x"779", x"77a", x"77b", x"77d", x"77e", 
    x"77f", x"780", x"781", x"782", x"783", x"784", x"785", x"786", 
    x"787", x"788", x"789", x"78a", x"78c", x"78d", x"78e", x"78f", 
    x"790", x"791", x"792", x"793", x"794", x"795", x"796", x"797", 
    x"798", x"799", x"79a", x"79b", x"79c", x"79d", x"79e", x"79e", 
    x"79f", x"7a0", x"7a1", x"7a2", x"7a3", x"7a4", x"7a5", x"7a6", 
    x"7a7", x"7a8", x"7a9", x"7aa", x"7aa", x"7ab", x"7ac", x"7ad", 
    x"7ae", x"7af", x"7b0", x"7b1", x"7b1", x"7b2", x"7b3", x"7b4", 
    x"7b5", x"7b6", x"7b7", x"7b7", x"7b8", x"7b9", x"7ba", x"7bb", 
    x"7bb", x"7bc", x"7bd", x"7be", x"7bf", x"7bf", x"7c0", x"7c1", 
    x"7c2", x"7c2", x"7c3", x"7c4", x"7c5", x"7c5", x"7c6", x"7c7", 
    x"7c8", x"7c8", x"7c9", x"7ca", x"7ca", x"7cb", x"7cc", x"7cd", 
    x"7cd", x"7ce", x"7cf", x"7cf", x"7d0", x"7d1", x"7d1", x"7d2", 
    x"7d3", x"7d3", x"7d4", x"7d5", x"7d5", x"7d6", x"7d6", x"7d7", 
    x"7d8", x"7d8", x"7d9", x"7d9", x"7da", x"7db", x"7db", x"7dc", 
    x"7dc", x"7dd", x"7de", x"7de", x"7df", x"7df", x"7e0", x"7e0", 
    x"7e1", x"7e1", x"7e2", x"7e2", x"7e3", x"7e3", x"7e4", x"7e5", 
    x"7e5", x"7e6", x"7e6", x"7e6", x"7e7", x"7e7", x"7e8", x"7e8", 
    x"7e9", x"7e9", x"7ea", x"7ea", x"7eb", x"7eb", x"7ec", x"7ec", 
    x"7ec", x"7ed", x"7ed", x"7ee", x"7ee", x"7ee", x"7ef", x"7ef", 
    x"7f0", x"7f0", x"7f0", x"7f1", x"7f1", x"7f1", x"7f2", x"7f2", 
    x"7f3", x"7f3", x"7f3", x"7f4", x"7f4", x"7f4", x"7f5", x"7f5", 
    x"7f5", x"7f5", x"7f6", x"7f6", x"7f6", x"7f7", x"7f7", x"7f7", 
    x"7f7", x"7f8", x"7f8", x"7f8", x"7f8", x"7f9", x"7f9", x"7f9", 
    x"7f9", x"7fa", x"7fa", x"7fa", x"7fa", x"7fb", x"7fb", x"7fb", 
    x"7fb", x"7fb", x"7fc", x"7fc", x"7fc", x"7fc", x"7fc", x"7fc", 
    x"7fd", x"7fd", x"7fd", x"7fd", x"7fd", x"7fd", x"7fd", x"7fd", 
    x"7fe", x"7fe", x"7fe", x"7fe", x"7fe", x"7fe", x"7fe", x"7fe", 
    x"7fe", x"7fe", x"7ff", x"7ff", x"7ff", x"7ff", x"7ff", x"7ff", 
    x"7ff", x"7ff", x"7ff", x"7ff", x"7ff", x"7ff", x"7ff", x"7ff");


begin

PROCESS (CLK)
BEGIN
	if (rising_edge (clk)) then
		sin <= isin(conv_integer(ADD));
		cos <= icos(conv_integer(ADD));		
	end if;
END PROCESS;


end architecture;
