software/prom-generic-dp-32.vhd