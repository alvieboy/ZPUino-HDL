library IEEE;
use IEEE.std_logic_1164.all; 
use IEEE.std_logic_unsigned.all; 
use ieee.numeric_std.all;

entity bootloader_dp_32 is
  port (
    CLK:              in std_logic;
    WEA:  in std_logic;
    ENA:  in std_logic;
    MASKA:    in std_logic_vector(3 downto 0);
    ADDRA:         in std_logic_vector(11 downto 2);
    DIA:        in std_logic_vector(31 downto 0);
    DOA:         out std_logic_vector(31 downto 0);
    WEB:  in std_logic;
    ENB:  in std_logic;
    ADDRB:         in std_logic_vector(11 downto 2);
    DIB:        in std_logic_vector(31 downto 0);
    MASKB:    in std_logic_vector(3 downto 0);
    DOB:         out std_logic_vector(31 downto 0)
  );
end entity bootloader_dp_32;

architecture behave of bootloader_dp_32 is

  subtype RAM_WORD is STD_LOGIC_VECTOR (31 downto 0);
  type RAM_TABLE is array (0 to 1023) of RAM_WORD;
 shared variable RAM: RAM_TABLE := RAM_TABLE'(
x"0b0b0b99",x"bf040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b99",x"9d040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fd0608",x"72830609",x"81058205",x"832b2a83",x"ffff0652",x"04000000",x"00000000",x"00000000",x"71fd0608",x"83ffff73",x"83060981",x"05820583",x"2b2b0906",x"7383ffff",x"0b0b0b0b",x"83a70400",x"72098105",x"72057373",x"09060906",x"73097306",x"070a8106",x"53510400",x"00000000",x"00000000",x"72722473",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71737109",x"71068106",x"30720a10",x"0a720a10",x"0a31050a",x"81065151",x"53510400",x"00000000",x"72722673",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"cc040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"720a722b",x"0a535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72729f06",x"0981050b",x"0b0b88af",x"05040000",x"00000000",x"00000000",x"00000000",x"00000000",x"72722aff",x"739f062a",x"0974090a",x"8106ff05",x"06075351",x"04000000",x"00000000",x"00000000",x"71715351",x"020d0406",x"73830609",x"81058205",x"832b0b2b",x"0772fc06",x"0c515104",x"00000000",x"72098105",x"72050970",x"81050906",x"0a810653",x"51040000",x"00000000",x"00000000",x"00000000",x"72098105",x"72050970",x"81050906",x"0a098106",x"53510400",x"00000000",x"00000000",x"00000000",x"71098105",x"52040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72720981",x"05055351",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097206",x"73730906",x"07535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fc0608",x"72830609",x"81058305",x"1010102a",x"81ff0652",x"04000000",x"00000000",x"00000000",x"71fc0608",x"0b0b0b9c",x"cc738306",x"10100508",x"060b0b0b",x"88b20400",x"00000000",x"00000000",x"0b0b0b89",x"80040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"e8040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097081",x"0509060a",x"8106ff05",x"70547106",x"73097274",x"05ff0506",x"07515151",x"04000000",x"72097081",x"0509060a",x"098106ff",x"05705471",x"06730972",x"7405ff05",x"06075151",x"51040000",x"05ff0504",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"810b0b0b",x"0b9d840c",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71810552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"02840572",x"10100552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"717105ff",x"05715351",x"020d0400",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"81dd3f94",x"9d3f0400",x"00000000",x"00000000",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101053",x"51047381",x"ff067383",x"06098105",x"83051010",x"102b0772",x"fc060c51",x"51043c04",x"72728072",x"8106ff05",x"09720605",x"71105272",x"0a100a53",x"72ed3851",x"51535104",x"88088c08",x"90087575",x"9b8d2d50",x"50880856",x"900c8c0c",x"880c5104",x"88088c08",x"90087575",x"9ac92d50",x"50880856",x"900c8c0c",x"880c5104",x"88088c08",x"90088eea",x"2d900c8c",x"0c880c04",x"ff3d0d0b",x"0b0b9da8",x"335170a6",x"389d9008",x"70085252",x"70802e92",x"3884129d",x"900c702d",x"9d900870",x"08525270",x"f038810b",x"0b0b0b9d",x"a834833d",x"0d040480",x"3d0d0b0b",x"0b9dd408",x"802e8e38",x"0b0b0b0b",x"800b802e",x"09810685",x"38823d0d",x"040b0b0b",x"9dd4510b",x"0b0bf5f8",x"3f823d0d",x"0404ff3d",x"0d80c480",x"80845271",x"0870822a",x"70810651",x"515170f3",x"38833d0d",x"04ff3d0d",x"80c48080",x"84527108",x"70812a70",x"81065151",x"5170f338",x"7382900a",x"0c833d0d",x"04ff3d0d",x"80c48080",x"84527108",x"70812a70",x"81065151",x"5170f338",x"7382900a",x"0c833d0d",x"04ff3d0d",x"738f0652",x"89722787",x"3880d712",x"518439b0",x"12518ac9",x"2d833d0d",x"04ff3d0d",x"7370842a",x"52528ae9",x"2d71518a",x"e92d833d",x"0d04ff3d",x"0d737098",x"2a52528b",x"852d7190",x"2a518b85",x"2d71882a",x"518b852d",x"71518b85",x"2d833d0d",x"04fe3d0d",x"747080dc",x"8080880c",x"7081ff06",x"ff831154",x"51537181",x"268d3880",x"fd518ac9",x"2d72a032",x"51833972",x"518ac92d",x"843d0d04",x"803d0d83",x"ffff0b83",x"d00a0c80",x"fe518ac9",x"2d823d0d",x"04ff3d0d",x"83d00a08",x"70882a52",x"528bbd2d",x"7181ff06",x"518bbd2d",x"80fe518a",x"c92d833d",x"0d0482f6",x"ff0b80cc",x"8080880c",x"800b80cc",x"8080840c",x"9f0b8390",x"0a0c04ff",x"3d0d7370",x"08515180",x"c8808084",x"70087084",x"80800772",x"0c525283",x"3d0d04ff",x"3d0d80c8",x"80808470",x"0870fbff",x"ff06720c",x"5252833d",x"0d04a090",x"0ba0800c",x"9dac0ba0",x"840c9995",x"2dff3d0d",x"73518b71",x"0c901152",x"98808072",x"0c80720c",x"700883ff",x"ff06880c",x"833d0d04",x"fa3d0d78",x"7a7dff1e",x"57575853",x"73ff2ea7",x"38805684",x"5275730c",x"72088818",x"0cff1252",x"71f33874",x"84167408",x"720cff16",x"56565273",x"ff2e0981",x"06dd3888",x"3d0d04f9",x"3d0d80d0",x"80808456",x"83d00a58",x"8cd72d75",x"518cfd2d",x"9dac7088",x"08101098",x"80840571",x"70840553",x"0c5657fb",x"8084a1ad",x"750c9d94",x"0b88180c",x"8070770c",x"760c7508",x"7083ffff",x"06515783",x"ffff780c",x"a0805488",x"08537752",x"75518d9c",x"2d75518c",x"bb2d7708",x"5574772e",x"893880c3",x"518ac92d",x"ff39a084",x"085574fb",x"a090ae80",x"2e893880",x"c2518ac9",x"2dff3980",x"d00a7008",x"70ffbf06",x"720c5656",x"8a8e2d8c",x"ee2dff3d",x"0d9db808",x"81119db8",x"0c518390",x"0a700870",x"feff0672",x"0c525283",x"3d0d0480",x"3d0d8bec",x"2d728180",x"07518bbd",x"2d8c812d",x"823d0d04",x"fe3d0d80",x"d0808084",x"538cd72d",x"85730c80",x"730c7208",x"7081ff06",x"74535152",x"8cbb2d71",x"880c843d",x"0d04fc3d",x"0d768111",x"33821233",x"7181800a",x"29718480",x"80290583",x"14337082",x"80291284",x"16335271",x"05a08005",x"86168517",x"33575253",x"53555755",x"53ff1353",x"72ff2e91",x"38737081",x"05553352",x"71757081",x"055734e9",x"3989518f",x"872d863d",x"0d04f93d",x"0d795780",x"d0808084",x"568cd72d",x"81173382",x"18337182",x"80290553",x"5371802e",x"94388517",x"72555372",x"70810554",x"33760cff",x"145473f3",x"38831733",x"84183371",x"82802905",x"56528054",x"73752797",x"38735877",x"760c7317",x"76085353",x"71733481",x"14547474",x"26ed3875",x"518cbb2d",x"8bec2d81",x"84518bbd",x"2d74882a",x"518bbd2d",x"74518bbd",x"2d805473",x"75278f38",x"73177033",x"52528bbd",x"2d811454",x"ee398c81",x"2d893d0d",x"04f93d0d",x"795680d0",x"80808455",x"8cd72d86",x"750c7451",x"8cbb2d8c",x"d72d81ad",x"70760c81",x"17338218",x"33718280",x"29058319",x"33780c84",x"1933780c",x"85193378",x"0c595353",x"80547377",x"27b33872",x"5873802e",x"87388cd7",x"2d77750c",x"73168611",x"33760c87",x"1133760c",x"5274518c",x"bb2d8f9c",x"2d880881",x"065271f6",x"38821454",x"767426d1",x"388cd72d",x"84750c74",x"518cbb2d",x"8bec2d81",x"87518bbd",x"2d8c812d",x"893d0d04",x"fc3d0d76",x"81113382",x"12337190",x"2b71882b",x"07831433",x"70720788",x"2b841633",x"71075152",x"53575754",x"5288518f",x"872d81ff",x"518ac92d",x"80c48080",x"84537208",x"70812a70",x"81065151",x"5271f338",x"73848080",x"0780c480",x"80840c86",x"3d0d04fe",x"3d0d8f9c",x"2d880888",x"08810653",x"5371f338",x"8bec2d81",x"83518bbd",x"2d72518b",x"bd2d8c81",x"2d843d0d",x"04fe3d0d",x"800b9db8",x"0c8bec2d",x"8181518b",x"bd2d9d94",x"53935272",x"70810554",x"33518bbd",x"2dff1252",x"71ff2e09",x"8106ec38",x"8c812d84",x"3d0d04fe",x"3d0d800b",x"9db80c8b",x"ec2d8182",x"518bbd2d",x"80d08080",x"84528cd7",x"2d81f90a",x"0b80d080",x"809c0c71",x"08725253",x"8cbb2d72",x"9dc00c72",x"902a518b",x"bd2d9dc0",x"08882a51",x"8bbd2d9d",x"c008518b",x"bd2d8f9c",x"2d880851",x"8bbd2d8c",x"812d843d",x"0d04803d",x"0d810b9d",x"bc0c800b",x"83900a0c",x"85518f87",x"2d823d0d",x"04803d0d",x"800b9dbc",x"0c8ca22d",x"86518f87",x"2d823d0d",x"04fd3d0d",x"80d08080",x"84548a51",x"8f872d8c",x"d72d9dac",x"7452538c",x"fd2d7288",x"08101098",x"80840571",x"70840553",x"0c52fb80",x"84a1ad72",x"0c9d940b",x"88140c73",x"518cbb2d",x"8a8e2d8c",x"ee2d8480",x"b30b80c4",x"8080840c",x"04ffab3d",x"0d80d93d",x"0856800b",x"9dbc0c80",x"0b9db80c",x"800bdf80",x"179d9971",x"902a7156",x"56575557",x"72727081",x"05543473",x"882a5372",x"72347382",x"16347598",x"2a52718b",x"16347590",x"2a52718c",x"16347588",x"2a52718d",x"1634758e",x"16348eea",x"0ba0800c",x"80c48080",x"84558480",x"b3750c80",x"c88080a4",x"53fbffff",x"73087072",x"06750c53",x"5480c880",x"80947008",x"70760672",x"0c535388",x"0b80c080",x"80840c90",x"0a538173",x"0c8ca22d",x"fe88880b",x"80dc8080",x"840c81f2",x"0b80d00a",x"0c80d080",x"80847052",x"528cbb2d",x"8cd72d71",x"518cbb2d",x"8cd72d84",x"720c7151",x"8cbb2d76",x"77767593",x"3d41415b",x"5b5b83d0",x"0a5c7808",x"70810651",x"52719d38",x"9dbc0853",x"72f0389d",x"b8085287",x"e87227e6",x"38727e0c",x"7283900a",x"0c998d2d",x"82900a08",x"5379802e",x"81b43872",x"80fe2e09",x"810680f4",x"3876802e",x"c138807d",x"7857575a",x"827727ff",x"b53883ff",x"ff7c0c79",x"fe185353",x"79722798",x"3880dc80",x"80887255",x"58721670",x"33790c52",x"81135373",x"7326f238",x"ff157611",x"547605ff",x"05703374",x"33707288",x"2b077f08",x"53515551",x"5271732e",x"098106fe",x"ed387533",x"53728a26",x"fee43872",x"10109cd8",x"05765270",x"08515271",x"2dfed339",x"7280fd2e",x"09810686",x"38815bfe",x"c5397682",x"9f269e38",x"7a802e87",x"388073a0",x"32545b80",x"d73d7705",x"fde00552",x"72723481",x"1757fea2",x"39805afe",x"9d397280",x"fe2e0981",x"06fe9338",x"7957ff7c",x"0c81775c",x"5afe8739",x"ff3d0d9a",x"9d2d7352",x"805195b1",x"2d833d0d",x"0483ffff",x"f80d8dd7",x"0483ffff",x"f80da088",x"04880880",x"c0808088",x"08a08008",x"2d50880c",x"810b900a",x"0c048d0b",x"8aa92d50",x"8a0b8aa9",x"2d500495",x"a62dbe0b",x"8aa92d50",x"99b22d80",x"700cfaad",x"95b4da0b",x"81808070",x"8b9a2d50",x"ad0b8aa9",x"2d50718b",x"9a2d5071",x"710c7180",x"08bd0b8a",x"a92d5070",x"0b8b9a2d",x"5099b22d",x"2e873870",x"115199d7",x"045198fc",x"2d000000",x"00000000",x"820b80c0",x"8080900c",x"0b0b0b04",x"0083f00a",x"0b800ba0",x"80721208",x"720c8412",x"5271712e",x"ff05f238",x"028c050d",x"9a900400",x"00000000",x"00000000",x"00000000",x"00fb3d0d",x"77795555",x"80567575",x"24ab3880",x"74249d38",x"80537352",x"745180e1",x"3f880854",x"75802e85",x"38880830",x"5473880c",x"873d0d04",x"73307681",x"325754dc",x"39743055",x"81567380",x"25d238ec",x"39fa3d0d",x"787a5755",x"80577675",x"24a43875",x"9f2c5481",x"53757432",x"74315274",x"519b3f88",x"08547680",x"2e853888",x"08305473",x"880c883d",x"0d047430",x"558157d7",x"39fc3d0d",x"76785354",x"81538074",x"73265255",x"72802e98",x"3870802e",x"a9388072",x"24a43871",x"10731075",x"72265354",x"5272ea38",x"73517883",x"38745170",x"880c863d",x"0d047281",x"2a72812a",x"53537280",x"2ee63871",x"7426ef38",x"73723175",x"74077481",x"2a74812a",x"55555654",x"e539ff3d",x"0d9dc80b",x"fc057008",x"525270ff",x"2e913870",x"2dfc1270",x"08525270",x"ff2e0981",x"06f13883",x"3d0d0404",x"ecde3f04",x"00ffffff",x"ff00ffff",x"ffff00ff",x"ffffff00",x"000009b1",x"000009e3",x"0000098b",x"00000816",x"00000a3a",x"00000a51",x"000008a9",x"00000938",x"000007c2",x"00000a65",x"00000000",x"00000000",x"00000000",x"00000ed0",x"01090600",x"00000000",x"05b8d800",x"b4041700",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"ffffffff",x"00000000",x"ffffffff",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000");

begin

  process (clk)
  begin
    if rising_edge(clk) then
      if ENA='1' then
        if WEA='1' then
          RAM(conv_integer(ADDRA) ) := DIA;
        end if;
        DOA <= RAM(conv_integer(ADDRA)) ;
      end if;
    end if;
  end process;  

  process (clk)
  begin
    if rising_edge(clk) then
      if ENB='1' then
        if WEB='1' then
          RAM( conv_integer(ADDRB) ) := DIB;
        end if;
        DOB <= RAM(conv_integer(ADDRB)) ;
      end if;
    end if;
  end process;  
end behave;
