bootloader/prom-generic-dp-32.vhd