---------------------------------------------------------------------
--	Filename:	gh_nsincos_rom_16_4.vhd
--			
--	Description:
--		- Sin Cos look up table 16 bit (from 1/4 table)
--
--	Copyright (c) 2008, 2009 by George Huber 
--		an OpenCores.org Project
--		free to use, but see documentation for conditions 
--
--	Revision 	History:
--	Revision 	Date      	Author   	Comment
--	-------- 	----------	---------	-----------
--	1.0      	11/01/08  	h LeFevre	Initial revision
--	2.0     	03/07/09  	h LeFevre	correct port name
--	
------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.STD_LOGIC_arith.all;
use IEEE.std_logic_unsigned.all;

entity gh_nsincos_rom_16_4 is
	port (
		CLK : in std_logic;
		ADD : in std_logic_vector(15 downto 0);
		nsin : out std_logic_vector(15 downto 0);
		cos : out std_logic_vector(15 downto 0)
		);
end entity;

architecture a of gh_nsincos_rom_16_4 is

	signal pdsADD, pdcADD :  STD_LOGIC;
	signal dsADD, dcADD :  STD_LOGIC;
	signal sAz, cAz   :  STD_LOGIC;
	signal sADD, cADD :  STD_LOGIC_VECTOR(15 DOWNTO 0);
	signal msin, mcos :  STD_LOGIC_VECTOR(15 DOWNTO 0);

	type rom_mem is array (0 to 16383) of std_logic_vector (15 downto 0);
	constant isin : rom_mem :=(  
    x"0000", x"0003", x"0006", x"0009", x"000d", x"0010", x"0013", x"0016", 
    x"0019", x"001c", x"001f", x"0023", x"0026", x"0029", x"002c", x"002f", 
    x"0032", x"0035", x"0039", x"003c", x"003f", x"0042", x"0045", x"0048", 
    x"004b", x"004f", x"0052", x"0055", x"0058", x"005b", x"005e", x"0061", 
    x"0065", x"0068", x"006b", x"006e", x"0071", x"0074", x"0077", x"007b", 
    x"007e", x"0081", x"0084", x"0087", x"008a", x"008d", x"0091", x"0094", 
    x"0097", x"009a", x"009d", x"00a0", x"00a3", x"00a6", x"00aa", x"00ad", 
    x"00b0", x"00b3", x"00b6", x"00b9", x"00bc", x"00c0", x"00c3", x"00c6", 
    x"00c9", x"00cc", x"00cf", x"00d2", x"00d6", x"00d9", x"00dc", x"00df", 
    x"00e2", x"00e5", x"00e8", x"00ec", x"00ef", x"00f2", x"00f5", x"00f8", 
    x"00fb", x"00fe", x"0102", x"0105", x"0108", x"010b", x"010e", x"0111", 
    x"0114", x"0118", x"011b", x"011e", x"0121", x"0124", x"0127", x"012a", 
    x"012e", x"0131", x"0134", x"0137", x"013a", x"013d", x"0140", x"0144", 
    x"0147", x"014a", x"014d", x"0150", x"0153", x"0156", x"015a", x"015d", 
    x"0160", x"0163", x"0166", x"0169", x"016c", x"0170", x"0173", x"0176", 
    x"0179", x"017c", x"017f", x"0182", x"0186", x"0189", x"018c", x"018f", 
    x"0192", x"0195", x"0198", x"019c", x"019f", x"01a2", x"01a5", x"01a8", 
    x"01ab", x"01ae", x"01b2", x"01b5", x"01b8", x"01bb", x"01be", x"01c1", 
    x"01c4", x"01c8", x"01cb", x"01ce", x"01d1", x"01d4", x"01d7", x"01da", 
    x"01dd", x"01e1", x"01e4", x"01e7", x"01ea", x"01ed", x"01f0", x"01f3", 
    x"01f7", x"01fa", x"01fd", x"0200", x"0203", x"0206", x"0209", x"020d", 
    x"0210", x"0213", x"0216", x"0219", x"021c", x"021f", x"0223", x"0226", 
    x"0229", x"022c", x"022f", x"0232", x"0235", x"0239", x"023c", x"023f", 
    x"0242", x"0245", x"0248", x"024b", x"024f", x"0252", x"0255", x"0258", 
    x"025b", x"025e", x"0261", x"0265", x"0268", x"026b", x"026e", x"0271", 
    x"0274", x"0277", x"027b", x"027e", x"0281", x"0284", x"0287", x"028a", 
    x"028d", x"0291", x"0294", x"0297", x"029a", x"029d", x"02a0", x"02a3", 
    x"02a7", x"02aa", x"02ad", x"02b0", x"02b3", x"02b6", x"02b9", x"02bd", 
    x"02c0", x"02c3", x"02c6", x"02c9", x"02cc", x"02cf", x"02d2", x"02d6", 
    x"02d9", x"02dc", x"02df", x"02e2", x"02e5", x"02e8", x"02ec", x"02ef", 
    x"02f2", x"02f5", x"02f8", x"02fb", x"02fe", x"0302", x"0305", x"0308", 
    x"030b", x"030e", x"0311", x"0314", x"0318", x"031b", x"031e", x"0321", 
    x"0324", x"0327", x"032a", x"032e", x"0331", x"0334", x"0337", x"033a", 
    x"033d", x"0340", x"0344", x"0347", x"034a", x"034d", x"0350", x"0353", 
    x"0356", x"035a", x"035d", x"0360", x"0363", x"0366", x"0369", x"036c", 
    x"0370", x"0373", x"0376", x"0379", x"037c", x"037f", x"0382", x"0385", 
    x"0389", x"038c", x"038f", x"0392", x"0395", x"0398", x"039b", x"039f", 
    x"03a2", x"03a5", x"03a8", x"03ab", x"03ae", x"03b1", x"03b5", x"03b8", 
    x"03bb", x"03be", x"03c1", x"03c4", x"03c7", x"03cb", x"03ce", x"03d1", 
    x"03d4", x"03d7", x"03da", x"03dd", x"03e1", x"03e4", x"03e7", x"03ea", 
    x"03ed", x"03f0", x"03f3", x"03f7", x"03fa", x"03fd", x"0400", x"0403", 
    x"0406", x"0409", x"040d", x"0410", x"0413", x"0416", x"0419", x"041c", 
    x"041f", x"0423", x"0426", x"0429", x"042c", x"042f", x"0432", x"0435", 
    x"0438", x"043c", x"043f", x"0442", x"0445", x"0448", x"044b", x"044e", 
    x"0452", x"0455", x"0458", x"045b", x"045e", x"0461", x"0464", x"0468", 
    x"046b", x"046e", x"0471", x"0474", x"0477", x"047a", x"047e", x"0481", 
    x"0484", x"0487", x"048a", x"048d", x"0490", x"0494", x"0497", x"049a", 
    x"049d", x"04a0", x"04a3", x"04a6", x"04aa", x"04ad", x"04b0", x"04b3", 
    x"04b6", x"04b9", x"04bc", x"04bf", x"04c3", x"04c6", x"04c9", x"04cc", 
    x"04cf", x"04d2", x"04d5", x"04d9", x"04dc", x"04df", x"04e2", x"04e5", 
    x"04e8", x"04eb", x"04ef", x"04f2", x"04f5", x"04f8", x"04fb", x"04fe", 
    x"0501", x"0505", x"0508", x"050b", x"050e", x"0511", x"0514", x"0517", 
    x"051b", x"051e", x"0521", x"0524", x"0527", x"052a", x"052d", x"0530", 
    x"0534", x"0537", x"053a", x"053d", x"0540", x"0543", x"0546", x"054a", 
    x"054d", x"0550", x"0553", x"0556", x"0559", x"055c", x"0560", x"0563", 
    x"0566", x"0569", x"056c", x"056f", x"0572", x"0576", x"0579", x"057c", 
    x"057f", x"0582", x"0585", x"0588", x"058c", x"058f", x"0592", x"0595", 
    x"0598", x"059b", x"059e", x"05a1", x"05a5", x"05a8", x"05ab", x"05ae", 
    x"05b1", x"05b4", x"05b7", x"05bb", x"05be", x"05c1", x"05c4", x"05c7", 
    x"05ca", x"05cd", x"05d1", x"05d4", x"05d7", x"05da", x"05dd", x"05e0", 
    x"05e3", x"05e7", x"05ea", x"05ed", x"05f0", x"05f3", x"05f6", x"05f9", 
    x"05fc", x"0600", x"0603", x"0606", x"0609", x"060c", x"060f", x"0612", 
    x"0616", x"0619", x"061c", x"061f", x"0622", x"0625", x"0628", x"062c", 
    x"062f", x"0632", x"0635", x"0638", x"063b", x"063e", x"0642", x"0645", 
    x"0648", x"064b", x"064e", x"0651", x"0654", x"0657", x"065b", x"065e", 
    x"0661", x"0664", x"0667", x"066a", x"066d", x"0671", x"0674", x"0677", 
    x"067a", x"067d", x"0680", x"0683", x"0687", x"068a", x"068d", x"0690", 
    x"0693", x"0696", x"0699", x"069d", x"06a0", x"06a3", x"06a6", x"06a9", 
    x"06ac", x"06af", x"06b2", x"06b6", x"06b9", x"06bc", x"06bf", x"06c2", 
    x"06c5", x"06c8", x"06cc", x"06cf", x"06d2", x"06d5", x"06d8", x"06db", 
    x"06de", x"06e2", x"06e5", x"06e8", x"06eb", x"06ee", x"06f1", x"06f4", 
    x"06f7", x"06fb", x"06fe", x"0701", x"0704", x"0707", x"070a", x"070d", 
    x"0711", x"0714", x"0717", x"071a", x"071d", x"0720", x"0723", x"0727", 
    x"072a", x"072d", x"0730", x"0733", x"0736", x"0739", x"073c", x"0740", 
    x"0743", x"0746", x"0749", x"074c", x"074f", x"0752", x"0756", x"0759", 
    x"075c", x"075f", x"0762", x"0765", x"0768", x"076c", x"076f", x"0772", 
    x"0775", x"0778", x"077b", x"077e", x"0781", x"0785", x"0788", x"078b", 
    x"078e", x"0791", x"0794", x"0797", x"079b", x"079e", x"07a1", x"07a4", 
    x"07a7", x"07aa", x"07ad", x"07b1", x"07b4", x"07b7", x"07ba", x"07bd", 
    x"07c0", x"07c3", x"07c6", x"07ca", x"07cd", x"07d0", x"07d3", x"07d6", 
    x"07d9", x"07dc", x"07e0", x"07e3", x"07e6", x"07e9", x"07ec", x"07ef", 
    x"07f2", x"07f6", x"07f9", x"07fc", x"07ff", x"0802", x"0805", x"0808", 
    x"080b", x"080f", x"0812", x"0815", x"0818", x"081b", x"081e", x"0821", 
    x"0825", x"0828", x"082b", x"082e", x"0831", x"0834", x"0837", x"083a", 
    x"083e", x"0841", x"0844", x"0847", x"084a", x"084d", x"0850", x"0854", 
    x"0857", x"085a", x"085d", x"0860", x"0863", x"0866", x"086a", x"086d", 
    x"0870", x"0873", x"0876", x"0879", x"087c", x"087f", x"0883", x"0886", 
    x"0889", x"088c", x"088f", x"0892", x"0895", x"0899", x"089c", x"089f", 
    x"08a2", x"08a5", x"08a8", x"08ab", x"08ae", x"08b2", x"08b5", x"08b8", 
    x"08bb", x"08be", x"08c1", x"08c4", x"08c8", x"08cb", x"08ce", x"08d1", 
    x"08d4", x"08d7", x"08da", x"08dd", x"08e1", x"08e4", x"08e7", x"08ea", 
    x"08ed", x"08f0", x"08f3", x"08f7", x"08fa", x"08fd", x"0900", x"0903", 
    x"0906", x"0909", x"090c", x"0910", x"0913", x"0916", x"0919", x"091c", 
    x"091f", x"0922", x"0926", x"0929", x"092c", x"092f", x"0932", x"0935", 
    x"0938", x"093b", x"093f", x"0942", x"0945", x"0948", x"094b", x"094e", 
    x"0951", x"0955", x"0958", x"095b", x"095e", x"0961", x"0964", x"0967", 
    x"096a", x"096e", x"0971", x"0974", x"0977", x"097a", x"097d", x"0980", 
    x"0984", x"0987", x"098a", x"098d", x"0990", x"0993", x"0996", x"0999", 
    x"099d", x"09a0", x"09a3", x"09a6", x"09a9", x"09ac", x"09af", x"09b3", 
    x"09b6", x"09b9", x"09bc", x"09bf", x"09c2", x"09c5", x"09c8", x"09cc", 
    x"09cf", x"09d2", x"09d5", x"09d8", x"09db", x"09de", x"09e2", x"09e5", 
    x"09e8", x"09eb", x"09ee", x"09f1", x"09f4", x"09f7", x"09fb", x"09fe", 
    x"0a01", x"0a04", x"0a07", x"0a0a", x"0a0d", x"0a11", x"0a14", x"0a17", 
    x"0a1a", x"0a1d", x"0a20", x"0a23", x"0a26", x"0a2a", x"0a2d", x"0a30", 
    x"0a33", x"0a36", x"0a39", x"0a3c", x"0a3f", x"0a43", x"0a46", x"0a49", 
    x"0a4c", x"0a4f", x"0a52", x"0a55", x"0a59", x"0a5c", x"0a5f", x"0a62", 
    x"0a65", x"0a68", x"0a6b", x"0a6e", x"0a72", x"0a75", x"0a78", x"0a7b", 
    x"0a7e", x"0a81", x"0a84", x"0a87", x"0a8b", x"0a8e", x"0a91", x"0a94", 
    x"0a97", x"0a9a", x"0a9d", x"0aa1", x"0aa4", x"0aa7", x"0aaa", x"0aad", 
    x"0ab0", x"0ab3", x"0ab6", x"0aba", x"0abd", x"0ac0", x"0ac3", x"0ac6", 
    x"0ac9", x"0acc", x"0acf", x"0ad3", x"0ad6", x"0ad9", x"0adc", x"0adf", 
    x"0ae2", x"0ae5", x"0ae9", x"0aec", x"0aef", x"0af2", x"0af5", x"0af8", 
    x"0afb", x"0afe", x"0b02", x"0b05", x"0b08", x"0b0b", x"0b0e", x"0b11", 
    x"0b14", x"0b17", x"0b1b", x"0b1e", x"0b21", x"0b24", x"0b27", x"0b2a", 
    x"0b2d", x"0b31", x"0b34", x"0b37", x"0b3a", x"0b3d", x"0b40", x"0b43", 
    x"0b46", x"0b4a", x"0b4d", x"0b50", x"0b53", x"0b56", x"0b59", x"0b5c", 
    x"0b5f", x"0b63", x"0b66", x"0b69", x"0b6c", x"0b6f", x"0b72", x"0b75", 
    x"0b78", x"0b7c", x"0b7f", x"0b82", x"0b85", x"0b88", x"0b8b", x"0b8e", 
    x"0b92", x"0b95", x"0b98", x"0b9b", x"0b9e", x"0ba1", x"0ba4", x"0ba7", 
    x"0bab", x"0bae", x"0bb1", x"0bb4", x"0bb7", x"0bba", x"0bbd", x"0bc0", 
    x"0bc4", x"0bc7", x"0bca", x"0bcd", x"0bd0", x"0bd3", x"0bd6", x"0bd9", 
    x"0bdd", x"0be0", x"0be3", x"0be6", x"0be9", x"0bec", x"0bef", x"0bf3", 
    x"0bf6", x"0bf9", x"0bfc", x"0bff", x"0c02", x"0c05", x"0c08", x"0c0c", 
    x"0c0f", x"0c12", x"0c15", x"0c18", x"0c1b", x"0c1e", x"0c21", x"0c25", 
    x"0c28", x"0c2b", x"0c2e", x"0c31", x"0c34", x"0c37", x"0c3a", x"0c3e", 
    x"0c41", x"0c44", x"0c47", x"0c4a", x"0c4d", x"0c50", x"0c53", x"0c57", 
    x"0c5a", x"0c5d", x"0c60", x"0c63", x"0c66", x"0c69", x"0c6c", x"0c70", 
    x"0c73", x"0c76", x"0c79", x"0c7c", x"0c7f", x"0c82", x"0c85", x"0c89", 
    x"0c8c", x"0c8f", x"0c92", x"0c95", x"0c98", x"0c9b", x"0c9e", x"0ca2", 
    x"0ca5", x"0ca8", x"0cab", x"0cae", x"0cb1", x"0cb4", x"0cb7", x"0cbb", 
    x"0cbe", x"0cc1", x"0cc4", x"0cc7", x"0cca", x"0ccd", x"0cd1", x"0cd4", 
    x"0cd7", x"0cda", x"0cdd", x"0ce0", x"0ce3", x"0ce6", x"0cea", x"0ced", 
    x"0cf0", x"0cf3", x"0cf6", x"0cf9", x"0cfc", x"0cff", x"0d03", x"0d06", 
    x"0d09", x"0d0c", x"0d0f", x"0d12", x"0d15", x"0d18", x"0d1c", x"0d1f", 
    x"0d22", x"0d25", x"0d28", x"0d2b", x"0d2e", x"0d31", x"0d35", x"0d38", 
    x"0d3b", x"0d3e", x"0d41", x"0d44", x"0d47", x"0d4a", x"0d4e", x"0d51", 
    x"0d54", x"0d57", x"0d5a", x"0d5d", x"0d60", x"0d63", x"0d66", x"0d6a", 
    x"0d6d", x"0d70", x"0d73", x"0d76", x"0d79", x"0d7c", x"0d7f", x"0d83", 
    x"0d86", x"0d89", x"0d8c", x"0d8f", x"0d92", x"0d95", x"0d98", x"0d9c", 
    x"0d9f", x"0da2", x"0da5", x"0da8", x"0dab", x"0dae", x"0db1", x"0db5", 
    x"0db8", x"0dbb", x"0dbe", x"0dc1", x"0dc4", x"0dc7", x"0dca", x"0dce", 
    x"0dd1", x"0dd4", x"0dd7", x"0dda", x"0ddd", x"0de0", x"0de3", x"0de7", 
    x"0dea", x"0ded", x"0df0", x"0df3", x"0df6", x"0df9", x"0dfc", x"0e00", 
    x"0e03", x"0e06", x"0e09", x"0e0c", x"0e0f", x"0e12", x"0e15", x"0e19", 
    x"0e1c", x"0e1f", x"0e22", x"0e25", x"0e28", x"0e2b", x"0e2e", x"0e32", 
    x"0e35", x"0e38", x"0e3b", x"0e3e", x"0e41", x"0e44", x"0e47", x"0e4a", 
    x"0e4e", x"0e51", x"0e54", x"0e57", x"0e5a", x"0e5d", x"0e60", x"0e63", 
    x"0e67", x"0e6a", x"0e6d", x"0e70", x"0e73", x"0e76", x"0e79", x"0e7c", 
    x"0e80", x"0e83", x"0e86", x"0e89", x"0e8c", x"0e8f", x"0e92", x"0e95", 
    x"0e99", x"0e9c", x"0e9f", x"0ea2", x"0ea5", x"0ea8", x"0eab", x"0eae", 
    x"0eb1", x"0eb5", x"0eb8", x"0ebb", x"0ebe", x"0ec1", x"0ec4", x"0ec7", 
    x"0eca", x"0ece", x"0ed1", x"0ed4", x"0ed7", x"0eda", x"0edd", x"0ee0", 
    x"0ee3", x"0ee7", x"0eea", x"0eed", x"0ef0", x"0ef3", x"0ef6", x"0ef9", 
    x"0efc", x"0eff", x"0f03", x"0f06", x"0f09", x"0f0c", x"0f0f", x"0f12", 
    x"0f15", x"0f18", x"0f1c", x"0f1f", x"0f22", x"0f25", x"0f28", x"0f2b", 
    x"0f2e", x"0f31", x"0f35", x"0f38", x"0f3b", x"0f3e", x"0f41", x"0f44", 
    x"0f47", x"0f4a", x"0f4d", x"0f51", x"0f54", x"0f57", x"0f5a", x"0f5d", 
    x"0f60", x"0f63", x"0f66", x"0f6a", x"0f6d", x"0f70", x"0f73", x"0f76", 
    x"0f79", x"0f7c", x"0f7f", x"0f82", x"0f86", x"0f89", x"0f8c", x"0f8f", 
    x"0f92", x"0f95", x"0f98", x"0f9b", x"0f9f", x"0fa2", x"0fa5", x"0fa8", 
    x"0fab", x"0fae", x"0fb1", x"0fb4", x"0fb8", x"0fbb", x"0fbe", x"0fc1", 
    x"0fc4", x"0fc7", x"0fca", x"0fcd", x"0fd0", x"0fd4", x"0fd7", x"0fda", 
    x"0fdd", x"0fe0", x"0fe3", x"0fe6", x"0fe9", x"0fec", x"0ff0", x"0ff3", 
    x"0ff6", x"0ff9", x"0ffc", x"0fff", x"1002", x"1005", x"1009", x"100c", 
    x"100f", x"1012", x"1015", x"1018", x"101b", x"101e", x"1021", x"1025", 
    x"1028", x"102b", x"102e", x"1031", x"1034", x"1037", x"103a", x"103e", 
    x"1041", x"1044", x"1047", x"104a", x"104d", x"1050", x"1053", x"1056", 
    x"105a", x"105d", x"1060", x"1063", x"1066", x"1069", x"106c", x"106f", 
    x"1072", x"1076", x"1079", x"107c", x"107f", x"1082", x"1085", x"1088", 
    x"108b", x"108f", x"1092", x"1095", x"1098", x"109b", x"109e", x"10a1", 
    x"10a4", x"10a7", x"10ab", x"10ae", x"10b1", x"10b4", x"10b7", x"10ba", 
    x"10bd", x"10c0", x"10c3", x"10c7", x"10ca", x"10cd", x"10d0", x"10d3", 
    x"10d6", x"10d9", x"10dc", x"10e0", x"10e3", x"10e6", x"10e9", x"10ec", 
    x"10ef", x"10f2", x"10f5", x"10f8", x"10fc", x"10ff", x"1102", x"1105", 
    x"1108", x"110b", x"110e", x"1111", x"1114", x"1118", x"111b", x"111e", 
    x"1121", x"1124", x"1127", x"112a", x"112d", x"1130", x"1134", x"1137", 
    x"113a", x"113d", x"1140", x"1143", x"1146", x"1149", x"114c", x"1150", 
    x"1153", x"1156", x"1159", x"115c", x"115f", x"1162", x"1165", x"1168", 
    x"116c", x"116f", x"1172", x"1175", x"1178", x"117b", x"117e", x"1181", 
    x"1185", x"1188", x"118b", x"118e", x"1191", x"1194", x"1197", x"119a", 
    x"119d", x"11a1", x"11a4", x"11a7", x"11aa", x"11ad", x"11b0", x"11b3", 
    x"11b6", x"11b9", x"11bd", x"11c0", x"11c3", x"11c6", x"11c9", x"11cc", 
    x"11cf", x"11d2", x"11d5", x"11d9", x"11dc", x"11df", x"11e2", x"11e5", 
    x"11e8", x"11eb", x"11ee", x"11f1", x"11f5", x"11f8", x"11fb", x"11fe", 
    x"1201", x"1204", x"1207", x"120a", x"120d", x"1210", x"1214", x"1217", 
    x"121a", x"121d", x"1220", x"1223", x"1226", x"1229", x"122c", x"1230", 
    x"1233", x"1236", x"1239", x"123c", x"123f", x"1242", x"1245", x"1248", 
    x"124c", x"124f", x"1252", x"1255", x"1258", x"125b", x"125e", x"1261", 
    x"1264", x"1268", x"126b", x"126e", x"1271", x"1274", x"1277", x"127a", 
    x"127d", x"1280", x"1284", x"1287", x"128a", x"128d", x"1290", x"1293", 
    x"1296", x"1299", x"129c", x"12a0", x"12a3", x"12a6", x"12a9", x"12ac", 
    x"12af", x"12b2", x"12b5", x"12b8", x"12bb", x"12bf", x"12c2", x"12c5", 
    x"12c8", x"12cb", x"12ce", x"12d1", x"12d4", x"12d7", x"12db", x"12de", 
    x"12e1", x"12e4", x"12e7", x"12ea", x"12ed", x"12f0", x"12f3", x"12f7", 
    x"12fa", x"12fd", x"1300", x"1303", x"1306", x"1309", x"130c", x"130f", 
    x"1312", x"1316", x"1319", x"131c", x"131f", x"1322", x"1325", x"1328", 
    x"132b", x"132e", x"1332", x"1335", x"1338", x"133b", x"133e", x"1341", 
    x"1344", x"1347", x"134a", x"134d", x"1351", x"1354", x"1357", x"135a", 
    x"135d", x"1360", x"1363", x"1366", x"1369", x"136d", x"1370", x"1373", 
    x"1376", x"1379", x"137c", x"137f", x"1382", x"1385", x"1388", x"138c", 
    x"138f", x"1392", x"1395", x"1398", x"139b", x"139e", x"13a1", x"13a4", 
    x"13a8", x"13ab", x"13ae", x"13b1", x"13b4", x"13b7", x"13ba", x"13bd", 
    x"13c0", x"13c3", x"13c7", x"13ca", x"13cd", x"13d0", x"13d3", x"13d6", 
    x"13d9", x"13dc", x"13df", x"13e3", x"13e6", x"13e9", x"13ec", x"13ef", 
    x"13f2", x"13f5", x"13f8", x"13fb", x"13fe", x"1402", x"1405", x"1408", 
    x"140b", x"140e", x"1411", x"1414", x"1417", x"141a", x"141d", x"1421", 
    x"1424", x"1427", x"142a", x"142d", x"1430", x"1433", x"1436", x"1439", 
    x"143c", x"1440", x"1443", x"1446", x"1449", x"144c", x"144f", x"1452", 
    x"1455", x"1458", x"145c", x"145f", x"1462", x"1465", x"1468", x"146b", 
    x"146e", x"1471", x"1474", x"1477", x"147b", x"147e", x"1481", x"1484", 
    x"1487", x"148a", x"148d", x"1490", x"1493", x"1496", x"149a", x"149d", 
    x"14a0", x"14a3", x"14a6", x"14a9", x"14ac", x"14af", x"14b2", x"14b5", 
    x"14b9", x"14bc", x"14bf", x"14c2", x"14c5", x"14c8", x"14cb", x"14ce", 
    x"14d1", x"14d4", x"14d8", x"14db", x"14de", x"14e1", x"14e4", x"14e7", 
    x"14ea", x"14ed", x"14f0", x"14f3", x"14f7", x"14fa", x"14fd", x"1500", 
    x"1503", x"1506", x"1509", x"150c", x"150f", x"1512", x"1516", x"1519", 
    x"151c", x"151f", x"1522", x"1525", x"1528", x"152b", x"152e", x"1531", 
    x"1534", x"1538", x"153b", x"153e", x"1541", x"1544", x"1547", x"154a", 
    x"154d", x"1550", x"1553", x"1557", x"155a", x"155d", x"1560", x"1563", 
    x"1566", x"1569", x"156c", x"156f", x"1572", x"1576", x"1579", x"157c", 
    x"157f", x"1582", x"1585", x"1588", x"158b", x"158e", x"1591", x"1595", 
    x"1598", x"159b", x"159e", x"15a1", x"15a4", x"15a7", x"15aa", x"15ad", 
    x"15b0", x"15b3", x"15b7", x"15ba", x"15bd", x"15c0", x"15c3", x"15c6", 
    x"15c9", x"15cc", x"15cf", x"15d2", x"15d6", x"15d9", x"15dc", x"15df", 
    x"15e2", x"15e5", x"15e8", x"15eb", x"15ee", x"15f1", x"15f4", x"15f8", 
    x"15fb", x"15fe", x"1601", x"1604", x"1607", x"160a", x"160d", x"1610", 
    x"1613", x"1617", x"161a", x"161d", x"1620", x"1623", x"1626", x"1629", 
    x"162c", x"162f", x"1632", x"1635", x"1639", x"163c", x"163f", x"1642", 
    x"1645", x"1648", x"164b", x"164e", x"1651", x"1654", x"1657", x"165b", 
    x"165e", x"1661", x"1664", x"1667", x"166a", x"166d", x"1670", x"1673", 
    x"1676", x"167a", x"167d", x"1680", x"1683", x"1686", x"1689", x"168c", 
    x"168f", x"1692", x"1695", x"1698", x"169c", x"169f", x"16a2", x"16a5", 
    x"16a8", x"16ab", x"16ae", x"16b1", x"16b4", x"16b7", x"16ba", x"16be", 
    x"16c1", x"16c4", x"16c7", x"16ca", x"16cd", x"16d0", x"16d3", x"16d6", 
    x"16d9", x"16dc", x"16e0", x"16e3", x"16e6", x"16e9", x"16ec", x"16ef", 
    x"16f2", x"16f5", x"16f8", x"16fb", x"16fe", x"1702", x"1705", x"1708", 
    x"170b", x"170e", x"1711", x"1714", x"1717", x"171a", x"171d", x"1720", 
    x"1724", x"1727", x"172a", x"172d", x"1730", x"1733", x"1736", x"1739", 
    x"173c", x"173f", x"1742", x"1746", x"1749", x"174c", x"174f", x"1752", 
    x"1755", x"1758", x"175b", x"175e", x"1761", x"1764", x"1767", x"176b", 
    x"176e", x"1771", x"1774", x"1777", x"177a", x"177d", x"1780", x"1783", 
    x"1786", x"1789", x"178d", x"1790", x"1793", x"1796", x"1799", x"179c", 
    x"179f", x"17a2", x"17a5", x"17a8", x"17ab", x"17af", x"17b2", x"17b5", 
    x"17b8", x"17bb", x"17be", x"17c1", x"17c4", x"17c7", x"17ca", x"17cd", 
    x"17d0", x"17d4", x"17d7", x"17da", x"17dd", x"17e0", x"17e3", x"17e6", 
    x"17e9", x"17ec", x"17ef", x"17f2", x"17f6", x"17f9", x"17fc", x"17ff", 
    x"1802", x"1805", x"1808", x"180b", x"180e", x"1811", x"1814", x"1817", 
    x"181b", x"181e", x"1821", x"1824", x"1827", x"182a", x"182d", x"1830", 
    x"1833", x"1836", x"1839", x"183c", x"1840", x"1843", x"1846", x"1849", 
    x"184c", x"184f", x"1852", x"1855", x"1858", x"185b", x"185e", x"1861", 
    x"1865", x"1868", x"186b", x"186e", x"1871", x"1874", x"1877", x"187a", 
    x"187d", x"1880", x"1883", x"1886", x"188a", x"188d", x"1890", x"1893", 
    x"1896", x"1899", x"189c", x"189f", x"18a2", x"18a5", x"18a8", x"18ab", 
    x"18af", x"18b2", x"18b5", x"18b8", x"18bb", x"18be", x"18c1", x"18c4", 
    x"18c7", x"18ca", x"18cd", x"18d0", x"18d4", x"18d7", x"18da", x"18dd", 
    x"18e0", x"18e3", x"18e6", x"18e9", x"18ec", x"18ef", x"18f2", x"18f5", 
    x"18f9", x"18fc", x"18ff", x"1902", x"1905", x"1908", x"190b", x"190e", 
    x"1911", x"1914", x"1917", x"191a", x"191d", x"1921", x"1924", x"1927", 
    x"192a", x"192d", x"1930", x"1933", x"1936", x"1939", x"193c", x"193f", 
    x"1942", x"1946", x"1949", x"194c", x"194f", x"1952", x"1955", x"1958", 
    x"195b", x"195e", x"1961", x"1964", x"1967", x"196a", x"196e", x"1971", 
    x"1974", x"1977", x"197a", x"197d", x"1980", x"1983", x"1986", x"1989", 
    x"198c", x"198f", x"1993", x"1996", x"1999", x"199c", x"199f", x"19a2", 
    x"19a5", x"19a8", x"19ab", x"19ae", x"19b1", x"19b4", x"19b7", x"19bb", 
    x"19be", x"19c1", x"19c4", x"19c7", x"19ca", x"19cd", x"19d0", x"19d3", 
    x"19d6", x"19d9", x"19dc", x"19df", x"19e3", x"19e6", x"19e9", x"19ec", 
    x"19ef", x"19f2", x"19f5", x"19f8", x"19fb", x"19fe", x"1a01", x"1a04", 
    x"1a07", x"1a0b", x"1a0e", x"1a11", x"1a14", x"1a17", x"1a1a", x"1a1d", 
    x"1a20", x"1a23", x"1a26", x"1a29", x"1a2c", x"1a2f", x"1a32", x"1a36", 
    x"1a39", x"1a3c", x"1a3f", x"1a42", x"1a45", x"1a48", x"1a4b", x"1a4e", 
    x"1a51", x"1a54", x"1a57", x"1a5a", x"1a5e", x"1a61", x"1a64", x"1a67", 
    x"1a6a", x"1a6d", x"1a70", x"1a73", x"1a76", x"1a79", x"1a7c", x"1a7f", 
    x"1a82", x"1a85", x"1a89", x"1a8c", x"1a8f", x"1a92", x"1a95", x"1a98", 
    x"1a9b", x"1a9e", x"1aa1", x"1aa4", x"1aa7", x"1aaa", x"1aad", x"1ab1", 
    x"1ab4", x"1ab7", x"1aba", x"1abd", x"1ac0", x"1ac3", x"1ac6", x"1ac9", 
    x"1acc", x"1acf", x"1ad2", x"1ad5", x"1ad8", x"1adc", x"1adf", x"1ae2", 
    x"1ae5", x"1ae8", x"1aeb", x"1aee", x"1af1", x"1af4", x"1af7", x"1afa", 
    x"1afd", x"1b00", x"1b03", x"1b07", x"1b0a", x"1b0d", x"1b10", x"1b13", 
    x"1b16", x"1b19", x"1b1c", x"1b1f", x"1b22", x"1b25", x"1b28", x"1b2b", 
    x"1b2e", x"1b31", x"1b35", x"1b38", x"1b3b", x"1b3e", x"1b41", x"1b44", 
    x"1b47", x"1b4a", x"1b4d", x"1b50", x"1b53", x"1b56", x"1b59", x"1b5c", 
    x"1b60", x"1b63", x"1b66", x"1b69", x"1b6c", x"1b6f", x"1b72", x"1b75", 
    x"1b78", x"1b7b", x"1b7e", x"1b81", x"1b84", x"1b87", x"1b8a", x"1b8e", 
    x"1b91", x"1b94", x"1b97", x"1b9a", x"1b9d", x"1ba0", x"1ba3", x"1ba6", 
    x"1ba9", x"1bac", x"1baf", x"1bb2", x"1bb5", x"1bb9", x"1bbc", x"1bbf", 
    x"1bc2", x"1bc5", x"1bc8", x"1bcb", x"1bce", x"1bd1", x"1bd4", x"1bd7", 
    x"1bda", x"1bdd", x"1be0", x"1be3", x"1be7", x"1bea", x"1bed", x"1bf0", 
    x"1bf3", x"1bf6", x"1bf9", x"1bfc", x"1bff", x"1c02", x"1c05", x"1c08", 
    x"1c0b", x"1c0e", x"1c11", x"1c14", x"1c18", x"1c1b", x"1c1e", x"1c21", 
    x"1c24", x"1c27", x"1c2a", x"1c2d", x"1c30", x"1c33", x"1c36", x"1c39", 
    x"1c3c", x"1c3f", x"1c42", x"1c46", x"1c49", x"1c4c", x"1c4f", x"1c52", 
    x"1c55", x"1c58", x"1c5b", x"1c5e", x"1c61", x"1c64", x"1c67", x"1c6a", 
    x"1c6d", x"1c70", x"1c73", x"1c77", x"1c7a", x"1c7d", x"1c80", x"1c83", 
    x"1c86", x"1c89", x"1c8c", x"1c8f", x"1c92", x"1c95", x"1c98", x"1c9b", 
    x"1c9e", x"1ca1", x"1ca4", x"1ca8", x"1cab", x"1cae", x"1cb1", x"1cb4", 
    x"1cb7", x"1cba", x"1cbd", x"1cc0", x"1cc3", x"1cc6", x"1cc9", x"1ccc", 
    x"1ccf", x"1cd2", x"1cd5", x"1cd9", x"1cdc", x"1cdf", x"1ce2", x"1ce5", 
    x"1ce8", x"1ceb", x"1cee", x"1cf1", x"1cf4", x"1cf7", x"1cfa", x"1cfd", 
    x"1d00", x"1d03", x"1d06", x"1d09", x"1d0d", x"1d10", x"1d13", x"1d16", 
    x"1d19", x"1d1c", x"1d1f", x"1d22", x"1d25", x"1d28", x"1d2b", x"1d2e", 
    x"1d31", x"1d34", x"1d37", x"1d3a", x"1d3d", x"1d41", x"1d44", x"1d47", 
    x"1d4a", x"1d4d", x"1d50", x"1d53", x"1d56", x"1d59", x"1d5c", x"1d5f", 
    x"1d62", x"1d65", x"1d68", x"1d6b", x"1d6e", x"1d71", x"1d75", x"1d78", 
    x"1d7b", x"1d7e", x"1d81", x"1d84", x"1d87", x"1d8a", x"1d8d", x"1d90", 
    x"1d93", x"1d96", x"1d99", x"1d9c", x"1d9f", x"1da2", x"1da5", x"1da8", 
    x"1dac", x"1daf", x"1db2", x"1db5", x"1db8", x"1dbb", x"1dbe", x"1dc1", 
    x"1dc4", x"1dc7", x"1dca", x"1dcd", x"1dd0", x"1dd3", x"1dd6", x"1dd9", 
    x"1ddc", x"1ddf", x"1de3", x"1de6", x"1de9", x"1dec", x"1def", x"1df2", 
    x"1df5", x"1df8", x"1dfb", x"1dfe", x"1e01", x"1e04", x"1e07", x"1e0a", 
    x"1e0d", x"1e10", x"1e13", x"1e16", x"1e19", x"1e1d", x"1e20", x"1e23", 
    x"1e26", x"1e29", x"1e2c", x"1e2f", x"1e32", x"1e35", x"1e38", x"1e3b", 
    x"1e3e", x"1e41", x"1e44", x"1e47", x"1e4a", x"1e4d", x"1e50", x"1e54", 
    x"1e57", x"1e5a", x"1e5d", x"1e60", x"1e63", x"1e66", x"1e69", x"1e6c", 
    x"1e6f", x"1e72", x"1e75", x"1e78", x"1e7b", x"1e7e", x"1e81", x"1e84", 
    x"1e87", x"1e8a", x"1e8d", x"1e91", x"1e94", x"1e97", x"1e9a", x"1e9d", 
    x"1ea0", x"1ea3", x"1ea6", x"1ea9", x"1eac", x"1eaf", x"1eb2", x"1eb5", 
    x"1eb8", x"1ebb", x"1ebe", x"1ec1", x"1ec4", x"1ec7", x"1eca", x"1ece", 
    x"1ed1", x"1ed4", x"1ed7", x"1eda", x"1edd", x"1ee0", x"1ee3", x"1ee6", 
    x"1ee9", x"1eec", x"1eef", x"1ef2", x"1ef5", x"1ef8", x"1efb", x"1efe", 
    x"1f01", x"1f04", x"1f07", x"1f0a", x"1f0e", x"1f11", x"1f14", x"1f17", 
    x"1f1a", x"1f1d", x"1f20", x"1f23", x"1f26", x"1f29", x"1f2c", x"1f2f", 
    x"1f32", x"1f35", x"1f38", x"1f3b", x"1f3e", x"1f41", x"1f44", x"1f47", 
    x"1f4a", x"1f4e", x"1f51", x"1f54", x"1f57", x"1f5a", x"1f5d", x"1f60", 
    x"1f63", x"1f66", x"1f69", x"1f6c", x"1f6f", x"1f72", x"1f75", x"1f78", 
    x"1f7b", x"1f7e", x"1f81", x"1f84", x"1f87", x"1f8a", x"1f8d", x"1f91", 
    x"1f94", x"1f97", x"1f9a", x"1f9d", x"1fa0", x"1fa3", x"1fa6", x"1fa9", 
    x"1fac", x"1faf", x"1fb2", x"1fb5", x"1fb8", x"1fbb", x"1fbe", x"1fc1", 
    x"1fc4", x"1fc7", x"1fca", x"1fcd", x"1fd0", x"1fd3", x"1fd7", x"1fda", 
    x"1fdd", x"1fe0", x"1fe3", x"1fe6", x"1fe9", x"1fec", x"1fef", x"1ff2", 
    x"1ff5", x"1ff8", x"1ffb", x"1ffe", x"2001", x"2004", x"2007", x"200a", 
    x"200d", x"2010", x"2013", x"2016", x"2019", x"201c", x"2020", x"2023", 
    x"2026", x"2029", x"202c", x"202f", x"2032", x"2035", x"2038", x"203b", 
    x"203e", x"2041", x"2044", x"2047", x"204a", x"204d", x"2050", x"2053", 
    x"2056", x"2059", x"205c", x"205f", x"2062", x"2065", x"2068", x"206c", 
    x"206f", x"2072", x"2075", x"2078", x"207b", x"207e", x"2081", x"2084", 
    x"2087", x"208a", x"208d", x"2090", x"2093", x"2096", x"2099", x"209c", 
    x"209f", x"20a2", x"20a5", x"20a8", x"20ab", x"20ae", x"20b1", x"20b4", 
    x"20b7", x"20bb", x"20be", x"20c1", x"20c4", x"20c7", x"20ca", x"20cd", 
    x"20d0", x"20d3", x"20d6", x"20d9", x"20dc", x"20df", x"20e2", x"20e5", 
    x"20e8", x"20eb", x"20ee", x"20f1", x"20f4", x"20f7", x"20fa", x"20fd", 
    x"2100", x"2103", x"2106", x"2109", x"210c", x"2110", x"2113", x"2116", 
    x"2119", x"211c", x"211f", x"2122", x"2125", x"2128", x"212b", x"212e", 
    x"2131", x"2134", x"2137", x"213a", x"213d", x"2140", x"2143", x"2146", 
    x"2149", x"214c", x"214f", x"2152", x"2155", x"2158", x"215b", x"215e", 
    x"2161", x"2164", x"2168", x"216b", x"216e", x"2171", x"2174", x"2177", 
    x"217a", x"217d", x"2180", x"2183", x"2186", x"2189", x"218c", x"218f", 
    x"2192", x"2195", x"2198", x"219b", x"219e", x"21a1", x"21a4", x"21a7", 
    x"21aa", x"21ad", x"21b0", x"21b3", x"21b6", x"21b9", x"21bc", x"21bf", 
    x"21c2", x"21c5", x"21c9", x"21cc", x"21cf", x"21d2", x"21d5", x"21d8", 
    x"21db", x"21de", x"21e1", x"21e4", x"21e7", x"21ea", x"21ed", x"21f0", 
    x"21f3", x"21f6", x"21f9", x"21fc", x"21ff", x"2202", x"2205", x"2208", 
    x"220b", x"220e", x"2211", x"2214", x"2217", x"221a", x"221d", x"2220", 
    x"2223", x"2226", x"2229", x"222c", x"222f", x"2233", x"2236", x"2239", 
    x"223c", x"223f", x"2242", x"2245", x"2248", x"224b", x"224e", x"2251", 
    x"2254", x"2257", x"225a", x"225d", x"2260", x"2263", x"2266", x"2269", 
    x"226c", x"226f", x"2272", x"2275", x"2278", x"227b", x"227e", x"2281", 
    x"2284", x"2287", x"228a", x"228d", x"2290", x"2293", x"2296", x"2299", 
    x"229c", x"229f", x"22a2", x"22a5", x"22a9", x"22ac", x"22af", x"22b2", 
    x"22b5", x"22b8", x"22bb", x"22be", x"22c1", x"22c4", x"22c7", x"22ca", 
    x"22cd", x"22d0", x"22d3", x"22d6", x"22d9", x"22dc", x"22df", x"22e2", 
    x"22e5", x"22e8", x"22eb", x"22ee", x"22f1", x"22f4", x"22f7", x"22fa", 
    x"22fd", x"2300", x"2303", x"2306", x"2309", x"230c", x"230f", x"2312", 
    x"2315", x"2318", x"231b", x"231e", x"2321", x"2324", x"2327", x"232a", 
    x"232e", x"2331", x"2334", x"2337", x"233a", x"233d", x"2340", x"2343", 
    x"2346", x"2349", x"234c", x"234f", x"2352", x"2355", x"2358", x"235b", 
    x"235e", x"2361", x"2364", x"2367", x"236a", x"236d", x"2370", x"2373", 
    x"2376", x"2379", x"237c", x"237f", x"2382", x"2385", x"2388", x"238b", 
    x"238e", x"2391", x"2394", x"2397", x"239a", x"239d", x"23a0", x"23a3", 
    x"23a6", x"23a9", x"23ac", x"23af", x"23b2", x"23b5", x"23b8", x"23bb", 
    x"23be", x"23c1", x"23c4", x"23c7", x"23ca", x"23cd", x"23d0", x"23d4", 
    x"23d7", x"23da", x"23dd", x"23e0", x"23e3", x"23e6", x"23e9", x"23ec", 
    x"23ef", x"23f2", x"23f5", x"23f8", x"23fb", x"23fe", x"2401", x"2404", 
    x"2407", x"240a", x"240d", x"2410", x"2413", x"2416", x"2419", x"241c", 
    x"241f", x"2422", x"2425", x"2428", x"242b", x"242e", x"2431", x"2434", 
    x"2437", x"243a", x"243d", x"2440", x"2443", x"2446", x"2449", x"244c", 
    x"244f", x"2452", x"2455", x"2458", x"245b", x"245e", x"2461", x"2464", 
    x"2467", x"246a", x"246d", x"2470", x"2473", x"2476", x"2479", x"247c", 
    x"247f", x"2482", x"2485", x"2488", x"248b", x"248e", x"2491", x"2494", 
    x"2497", x"249a", x"249d", x"24a0", x"24a3", x"24a6", x"24a9", x"24ac", 
    x"24af", x"24b2", x"24b5", x"24b8", x"24bb", x"24be", x"24c1", x"24c5", 
    x"24c8", x"24cb", x"24ce", x"24d1", x"24d4", x"24d7", x"24da", x"24dd", 
    x"24e0", x"24e3", x"24e6", x"24e9", x"24ec", x"24ef", x"24f2", x"24f5", 
    x"24f8", x"24fb", x"24fe", x"2501", x"2504", x"2507", x"250a", x"250d", 
    x"2510", x"2513", x"2516", x"2519", x"251c", x"251f", x"2522", x"2525", 
    x"2528", x"252b", x"252e", x"2531", x"2534", x"2537", x"253a", x"253d", 
    x"2540", x"2543", x"2546", x"2549", x"254c", x"254f", x"2552", x"2555", 
    x"2558", x"255b", x"255e", x"2561", x"2564", x"2567", x"256a", x"256d", 
    x"2570", x"2573", x"2576", x"2579", x"257c", x"257f", x"2582", x"2585", 
    x"2588", x"258b", x"258e", x"2591", x"2594", x"2597", x"259a", x"259d", 
    x"25a0", x"25a3", x"25a6", x"25a9", x"25ac", x"25af", x"25b2", x"25b5", 
    x"25b8", x"25bb", x"25be", x"25c1", x"25c4", x"25c7", x"25ca", x"25cd", 
    x"25d0", x"25d3", x"25d6", x"25d9", x"25dc", x"25df", x"25e2", x"25e5", 
    x"25e8", x"25eb", x"25ee", x"25f1", x"25f4", x"25f7", x"25fa", x"25fd", 
    x"2600", x"2603", x"2606", x"2609", x"260c", x"260f", x"2612", x"2615", 
    x"2618", x"261b", x"261e", x"2621", x"2624", x"2627", x"262a", x"262d", 
    x"2630", x"2633", x"2636", x"2639", x"263c", x"263f", x"2642", x"2645", 
    x"2648", x"264b", x"264e", x"2651", x"2654", x"2657", x"265a", x"265d", 
    x"2660", x"2663", x"2666", x"2669", x"266c", x"266f", x"2672", x"2675", 
    x"2678", x"267b", x"267e", x"2681", x"2684", x"2687", x"268a", x"268d", 
    x"2690", x"2693", x"2696", x"2699", x"269c", x"269f", x"26a2", x"26a5", 
    x"26a8", x"26ab", x"26ae", x"26b1", x"26b4", x"26b7", x"26ba", x"26bd", 
    x"26c0", x"26c3", x"26c6", x"26c9", x"26cc", x"26cf", x"26d2", x"26d5", 
    x"26d8", x"26db", x"26de", x"26e1", x"26e4", x"26e7", x"26ea", x"26ed", 
    x"26f0", x"26f3", x"26f6", x"26f9", x"26fc", x"26ff", x"2702", x"2705", 
    x"2708", x"270b", x"270e", x"2711", x"2714", x"2717", x"271a", x"271d", 
    x"2720", x"2723", x"2726", x"2729", x"272c", x"272f", x"2731", x"2734", 
    x"2737", x"273a", x"273d", x"2740", x"2743", x"2746", x"2749", x"274c", 
    x"274f", x"2752", x"2755", x"2758", x"275b", x"275e", x"2761", x"2764", 
    x"2767", x"276a", x"276d", x"2770", x"2773", x"2776", x"2779", x"277c", 
    x"277f", x"2782", x"2785", x"2788", x"278b", x"278e", x"2791", x"2794", 
    x"2797", x"279a", x"279d", x"27a0", x"27a3", x"27a6", x"27a9", x"27ac", 
    x"27af", x"27b2", x"27b5", x"27b8", x"27bb", x"27be", x"27c1", x"27c4", 
    x"27c7", x"27ca", x"27cd", x"27d0", x"27d3", x"27d6", x"27d9", x"27dc", 
    x"27df", x"27e2", x"27e5", x"27e8", x"27eb", x"27ee", x"27f1", x"27f4", 
    x"27f7", x"27fa", x"27fd", x"2800", x"2803", x"2806", x"2809", x"280c", 
    x"280f", x"2812", x"2815", x"2817", x"281a", x"281d", x"2820", x"2823", 
    x"2826", x"2829", x"282c", x"282f", x"2832", x"2835", x"2838", x"283b", 
    x"283e", x"2841", x"2844", x"2847", x"284a", x"284d", x"2850", x"2853", 
    x"2856", x"2859", x"285c", x"285f", x"2862", x"2865", x"2868", x"286b", 
    x"286e", x"2871", x"2874", x"2877", x"287a", x"287d", x"2880", x"2883", 
    x"2886", x"2889", x"288c", x"288f", x"2892", x"2895", x"2898", x"289b", 
    x"289e", x"28a1", x"28a4", x"28a7", x"28aa", x"28ad", x"28b0", x"28b3", 
    x"28b5", x"28b8", x"28bb", x"28be", x"28c1", x"28c4", x"28c7", x"28ca", 
    x"28cd", x"28d0", x"28d3", x"28d6", x"28d9", x"28dc", x"28df", x"28e2", 
    x"28e5", x"28e8", x"28eb", x"28ee", x"28f1", x"28f4", x"28f7", x"28fa", 
    x"28fd", x"2900", x"2903", x"2906", x"2909", x"290c", x"290f", x"2912", 
    x"2915", x"2918", x"291b", x"291e", x"2921", x"2924", x"2927", x"292a", 
    x"292d", x"2930", x"2932", x"2935", x"2938", x"293b", x"293e", x"2941", 
    x"2944", x"2947", x"294a", x"294d", x"2950", x"2953", x"2956", x"2959", 
    x"295c", x"295f", x"2962", x"2965", x"2968", x"296b", x"296e", x"2971", 
    x"2974", x"2977", x"297a", x"297d", x"2980", x"2983", x"2986", x"2989", 
    x"298c", x"298f", x"2992", x"2995", x"2998", x"299b", x"299e", x"29a0", 
    x"29a3", x"29a6", x"29a9", x"29ac", x"29af", x"29b2", x"29b5", x"29b8", 
    x"29bb", x"29be", x"29c1", x"29c4", x"29c7", x"29ca", x"29cd", x"29d0", 
    x"29d3", x"29d6", x"29d9", x"29dc", x"29df", x"29e2", x"29e5", x"29e8", 
    x"29eb", x"29ee", x"29f1", x"29f4", x"29f7", x"29fa", x"29fd", x"29ff", 
    x"2a02", x"2a05", x"2a08", x"2a0b", x"2a0e", x"2a11", x"2a14", x"2a17", 
    x"2a1a", x"2a1d", x"2a20", x"2a23", x"2a26", x"2a29", x"2a2c", x"2a2f", 
    x"2a32", x"2a35", x"2a38", x"2a3b", x"2a3e", x"2a41", x"2a44", x"2a47", 
    x"2a4a", x"2a4d", x"2a50", x"2a53", x"2a56", x"2a58", x"2a5b", x"2a5e", 
    x"2a61", x"2a64", x"2a67", x"2a6a", x"2a6d", x"2a70", x"2a73", x"2a76", 
    x"2a79", x"2a7c", x"2a7f", x"2a82", x"2a85", x"2a88", x"2a8b", x"2a8e", 
    x"2a91", x"2a94", x"2a97", x"2a9a", x"2a9d", x"2aa0", x"2aa3", x"2aa6", 
    x"2aa8", x"2aab", x"2aae", x"2ab1", x"2ab4", x"2ab7", x"2aba", x"2abd", 
    x"2ac0", x"2ac3", x"2ac6", x"2ac9", x"2acc", x"2acf", x"2ad2", x"2ad5", 
    x"2ad8", x"2adb", x"2ade", x"2ae1", x"2ae4", x"2ae7", x"2aea", x"2aed", 
    x"2af0", x"2af2", x"2af5", x"2af8", x"2afb", x"2afe", x"2b01", x"2b04", 
    x"2b07", x"2b0a", x"2b0d", x"2b10", x"2b13", x"2b16", x"2b19", x"2b1c", 
    x"2b1f", x"2b22", x"2b25", x"2b28", x"2b2b", x"2b2e", x"2b31", x"2b34", 
    x"2b37", x"2b39", x"2b3c", x"2b3f", x"2b42", x"2b45", x"2b48", x"2b4b", 
    x"2b4e", x"2b51", x"2b54", x"2b57", x"2b5a", x"2b5d", x"2b60", x"2b63", 
    x"2b66", x"2b69", x"2b6c", x"2b6f", x"2b72", x"2b75", x"2b78", x"2b7b", 
    x"2b7d", x"2b80", x"2b83", x"2b86", x"2b89", x"2b8c", x"2b8f", x"2b92", 
    x"2b95", x"2b98", x"2b9b", x"2b9e", x"2ba1", x"2ba4", x"2ba7", x"2baa", 
    x"2bad", x"2bb0", x"2bb3", x"2bb6", x"2bb9", x"2bbb", x"2bbe", x"2bc1", 
    x"2bc4", x"2bc7", x"2bca", x"2bcd", x"2bd0", x"2bd3", x"2bd6", x"2bd9", 
    x"2bdc", x"2bdf", x"2be2", x"2be5", x"2be8", x"2beb", x"2bee", x"2bf1", 
    x"2bf4", x"2bf7", x"2bf9", x"2bfc", x"2bff", x"2c02", x"2c05", x"2c08", 
    x"2c0b", x"2c0e", x"2c11", x"2c14", x"2c17", x"2c1a", x"2c1d", x"2c20", 
    x"2c23", x"2c26", x"2c29", x"2c2c", x"2c2f", x"2c32", x"2c34", x"2c37", 
    x"2c3a", x"2c3d", x"2c40", x"2c43", x"2c46", x"2c49", x"2c4c", x"2c4f", 
    x"2c52", x"2c55", x"2c58", x"2c5b", x"2c5e", x"2c61", x"2c64", x"2c67", 
    x"2c6a", x"2c6c", x"2c6f", x"2c72", x"2c75", x"2c78", x"2c7b", x"2c7e", 
    x"2c81", x"2c84", x"2c87", x"2c8a", x"2c8d", x"2c90", x"2c93", x"2c96", 
    x"2c99", x"2c9c", x"2c9f", x"2ca1", x"2ca4", x"2ca7", x"2caa", x"2cad", 
    x"2cb0", x"2cb3", x"2cb6", x"2cb9", x"2cbc", x"2cbf", x"2cc2", x"2cc5", 
    x"2cc8", x"2ccb", x"2cce", x"2cd1", x"2cd4", x"2cd6", x"2cd9", x"2cdc", 
    x"2cdf", x"2ce2", x"2ce5", x"2ce8", x"2ceb", x"2cee", x"2cf1", x"2cf4", 
    x"2cf7", x"2cfa", x"2cfd", x"2d00", x"2d03", x"2d06", x"2d08", x"2d0b", 
    x"2d0e", x"2d11", x"2d14", x"2d17", x"2d1a", x"2d1d", x"2d20", x"2d23", 
    x"2d26", x"2d29", x"2d2c", x"2d2f", x"2d32", x"2d35", x"2d37", x"2d3a", 
    x"2d3d", x"2d40", x"2d43", x"2d46", x"2d49", x"2d4c", x"2d4f", x"2d52", 
    x"2d55", x"2d58", x"2d5b", x"2d5e", x"2d61", x"2d64", x"2d67", x"2d69", 
    x"2d6c", x"2d6f", x"2d72", x"2d75", x"2d78", x"2d7b", x"2d7e", x"2d81", 
    x"2d84", x"2d87", x"2d8a", x"2d8d", x"2d90", x"2d93", x"2d95", x"2d98", 
    x"2d9b", x"2d9e", x"2da1", x"2da4", x"2da7", x"2daa", x"2dad", x"2db0", 
    x"2db3", x"2db6", x"2db9", x"2dbc", x"2dbf", x"2dc2", x"2dc4", x"2dc7", 
    x"2dca", x"2dcd", x"2dd0", x"2dd3", x"2dd6", x"2dd9", x"2ddc", x"2ddf", 
    x"2de2", x"2de5", x"2de8", x"2deb", x"2dee", x"2df0", x"2df3", x"2df6", 
    x"2df9", x"2dfc", x"2dff", x"2e02", x"2e05", x"2e08", x"2e0b", x"2e0e", 
    x"2e11", x"2e14", x"2e17", x"2e19", x"2e1c", x"2e1f", x"2e22", x"2e25", 
    x"2e28", x"2e2b", x"2e2e", x"2e31", x"2e34", x"2e37", x"2e3a", x"2e3d", 
    x"2e40", x"2e42", x"2e45", x"2e48", x"2e4b", x"2e4e", x"2e51", x"2e54", 
    x"2e57", x"2e5a", x"2e5d", x"2e60", x"2e63", x"2e66", x"2e69", x"2e6b", 
    x"2e6e", x"2e71", x"2e74", x"2e77", x"2e7a", x"2e7d", x"2e80", x"2e83", 
    x"2e86", x"2e89", x"2e8c", x"2e8f", x"2e92", x"2e94", x"2e97", x"2e9a", 
    x"2e9d", x"2ea0", x"2ea3", x"2ea6", x"2ea9", x"2eac", x"2eaf", x"2eb2", 
    x"2eb5", x"2eb8", x"2eba", x"2ebd", x"2ec0", x"2ec3", x"2ec6", x"2ec9", 
    x"2ecc", x"2ecf", x"2ed2", x"2ed5", x"2ed8", x"2edb", x"2ede", x"2ee1", 
    x"2ee3", x"2ee6", x"2ee9", x"2eec", x"2eef", x"2ef2", x"2ef5", x"2ef8", 
    x"2efb", x"2efe", x"2f01", x"2f04", x"2f06", x"2f09", x"2f0c", x"2f0f", 
    x"2f12", x"2f15", x"2f18", x"2f1b", x"2f1e", x"2f21", x"2f24", x"2f27", 
    x"2f2a", x"2f2c", x"2f2f", x"2f32", x"2f35", x"2f38", x"2f3b", x"2f3e", 
    x"2f41", x"2f44", x"2f47", x"2f4a", x"2f4d", x"2f50", x"2f52", x"2f55", 
    x"2f58", x"2f5b", x"2f5e", x"2f61", x"2f64", x"2f67", x"2f6a", x"2f6d", 
    x"2f70", x"2f73", x"2f75", x"2f78", x"2f7b", x"2f7e", x"2f81", x"2f84", 
    x"2f87", x"2f8a", x"2f8d", x"2f90", x"2f93", x"2f96", x"2f98", x"2f9b", 
    x"2f9e", x"2fa1", x"2fa4", x"2fa7", x"2faa", x"2fad", x"2fb0", x"2fb3", 
    x"2fb6", x"2fb9", x"2fbb", x"2fbe", x"2fc1", x"2fc4", x"2fc7", x"2fca", 
    x"2fcd", x"2fd0", x"2fd3", x"2fd6", x"2fd9", x"2fdb", x"2fde", x"2fe1", 
    x"2fe4", x"2fe7", x"2fea", x"2fed", x"2ff0", x"2ff3", x"2ff6", x"2ff9", 
    x"2ffc", x"2ffe", x"3001", x"3004", x"3007", x"300a", x"300d", x"3010", 
    x"3013", x"3016", x"3019", x"301c", x"301e", x"3021", x"3024", x"3027", 
    x"302a", x"302d", x"3030", x"3033", x"3036", x"3039", x"303c", x"303e", 
    x"3041", x"3044", x"3047", x"304a", x"304d", x"3050", x"3053", x"3056", 
    x"3059", x"305c", x"305e", x"3061", x"3064", x"3067", x"306a", x"306d", 
    x"3070", x"3073", x"3076", x"3079", x"307c", x"307e", x"3081", x"3084", 
    x"3087", x"308a", x"308d", x"3090", x"3093", x"3096", x"3099", x"309c", 
    x"309e", x"30a1", x"30a4", x"30a7", x"30aa", x"30ad", x"30b0", x"30b3", 
    x"30b6", x"30b9", x"30bc", x"30be", x"30c1", x"30c4", x"30c7", x"30ca", 
    x"30cd", x"30d0", x"30d3", x"30d6", x"30d9", x"30db", x"30de", x"30e1", 
    x"30e4", x"30e7", x"30ea", x"30ed", x"30f0", x"30f3", x"30f6", x"30f8", 
    x"30fb", x"30fe", x"3101", x"3104", x"3107", x"310a", x"310d", x"3110", 
    x"3113", x"3116", x"3118", x"311b", x"311e", x"3121", x"3124", x"3127", 
    x"312a", x"312d", x"3130", x"3133", x"3135", x"3138", x"313b", x"313e", 
    x"3141", x"3144", x"3147", x"314a", x"314d", x"3150", x"3152", x"3155", 
    x"3158", x"315b", x"315e", x"3161", x"3164", x"3167", x"316a", x"316c", 
    x"316f", x"3172", x"3175", x"3178", x"317b", x"317e", x"3181", x"3184", 
    x"3187", x"3189", x"318c", x"318f", x"3192", x"3195", x"3198", x"319b", 
    x"319e", x"31a1", x"31a4", x"31a6", x"31a9", x"31ac", x"31af", x"31b2", 
    x"31b5", x"31b8", x"31bb", x"31be", x"31c0", x"31c3", x"31c6", x"31c9", 
    x"31cc", x"31cf", x"31d2", x"31d5", x"31d8", x"31db", x"31dd", x"31e0", 
    x"31e3", x"31e6", x"31e9", x"31ec", x"31ef", x"31f2", x"31f5", x"31f7", 
    x"31fa", x"31fd", x"3200", x"3203", x"3206", x"3209", x"320c", x"320f", 
    x"3211", x"3214", x"3217", x"321a", x"321d", x"3220", x"3223", x"3226", 
    x"3229", x"322b", x"322e", x"3231", x"3234", x"3237", x"323a", x"323d", 
    x"3240", x"3243", x"3246", x"3248", x"324b", x"324e", x"3251", x"3254", 
    x"3257", x"325a", x"325d", x"325f", x"3262", x"3265", x"3268", x"326b", 
    x"326e", x"3271", x"3274", x"3277", x"3279", x"327c", x"327f", x"3282", 
    x"3285", x"3288", x"328b", x"328e", x"3291", x"3293", x"3296", x"3299", 
    x"329c", x"329f", x"32a2", x"32a5", x"32a8", x"32ab", x"32ad", x"32b0", 
    x"32b3", x"32b6", x"32b9", x"32bc", x"32bf", x"32c2", x"32c5", x"32c7", 
    x"32ca", x"32cd", x"32d0", x"32d3", x"32d6", x"32d9", x"32dc", x"32de", 
    x"32e1", x"32e4", x"32e7", x"32ea", x"32ed", x"32f0", x"32f3", x"32f6", 
    x"32f8", x"32fb", x"32fe", x"3301", x"3304", x"3307", x"330a", x"330d", 
    x"330f", x"3312", x"3315", x"3318", x"331b", x"331e", x"3321", x"3324", 
    x"3326", x"3329", x"332c", x"332f", x"3332", x"3335", x"3338", x"333b", 
    x"333e", x"3340", x"3343", x"3346", x"3349", x"334c", x"334f", x"3352", 
    x"3355", x"3357", x"335a", x"335d", x"3360", x"3363", x"3366", x"3369", 
    x"336c", x"336e", x"3371", x"3374", x"3377", x"337a", x"337d", x"3380", 
    x"3383", x"3385", x"3388", x"338b", x"338e", x"3391", x"3394", x"3397", 
    x"339a", x"339c", x"339f", x"33a2", x"33a5", x"33a8", x"33ab", x"33ae", 
    x"33b1", x"33b3", x"33b6", x"33b9", x"33bc", x"33bf", x"33c2", x"33c5", 
    x"33c8", x"33ca", x"33cd", x"33d0", x"33d3", x"33d6", x"33d9", x"33dc", 
    x"33df", x"33e1", x"33e4", x"33e7", x"33ea", x"33ed", x"33f0", x"33f3", 
    x"33f6", x"33f8", x"33fb", x"33fe", x"3401", x"3404", x"3407", x"340a", 
    x"340c", x"340f", x"3412", x"3415", x"3418", x"341b", x"341e", x"3421", 
    x"3423", x"3426", x"3429", x"342c", x"342f", x"3432", x"3435", x"3438", 
    x"343a", x"343d", x"3440", x"3443", x"3446", x"3449", x"344c", x"344e", 
    x"3451", x"3454", x"3457", x"345a", x"345d", x"3460", x"3463", x"3465", 
    x"3468", x"346b", x"346e", x"3471", x"3474", x"3477", x"3479", x"347c", 
    x"347f", x"3482", x"3485", x"3488", x"348b", x"348e", x"3490", x"3493", 
    x"3496", x"3499", x"349c", x"349f", x"34a2", x"34a4", x"34a7", x"34aa", 
    x"34ad", x"34b0", x"34b3", x"34b6", x"34b8", x"34bb", x"34be", x"34c1", 
    x"34c4", x"34c7", x"34ca", x"34cc", x"34cf", x"34d2", x"34d5", x"34d8", 
    x"34db", x"34de", x"34e1", x"34e3", x"34e6", x"34e9", x"34ec", x"34ef", 
    x"34f2", x"34f5", x"34f7", x"34fa", x"34fd", x"3500", x"3503", x"3506", 
    x"3509", x"350b", x"350e", x"3511", x"3514", x"3517", x"351a", x"351d", 
    x"351f", x"3522", x"3525", x"3528", x"352b", x"352e", x"3531", x"3533", 
    x"3536", x"3539", x"353c", x"353f", x"3542", x"3545", x"3547", x"354a", 
    x"354d", x"3550", x"3553", x"3556", x"3559", x"355b", x"355e", x"3561", 
    x"3564", x"3567", x"356a", x"356d", x"356f", x"3572", x"3575", x"3578", 
    x"357b", x"357e", x"3581", x"3583", x"3586", x"3589", x"358c", x"358f", 
    x"3592", x"3595", x"3597", x"359a", x"359d", x"35a0", x"35a3", x"35a6", 
    x"35a8", x"35ab", x"35ae", x"35b1", x"35b4", x"35b7", x"35ba", x"35bc", 
    x"35bf", x"35c2", x"35c5", x"35c8", x"35cb", x"35ce", x"35d0", x"35d3", 
    x"35d6", x"35d9", x"35dc", x"35df", x"35e1", x"35e4", x"35e7", x"35ea", 
    x"35ed", x"35f0", x"35f3", x"35f5", x"35f8", x"35fb", x"35fe", x"3601", 
    x"3604", x"3607", x"3609", x"360c", x"360f", x"3612", x"3615", x"3618", 
    x"361a", x"361d", x"3620", x"3623", x"3626", x"3629", x"362c", x"362e", 
    x"3631", x"3634", x"3637", x"363a", x"363d", x"363f", x"3642", x"3645", 
    x"3648", x"364b", x"364e", x"3651", x"3653", x"3656", x"3659", x"365c", 
    x"365f", x"3662", x"3664", x"3667", x"366a", x"366d", x"3670", x"3673", 
    x"3676", x"3678", x"367b", x"367e", x"3681", x"3684", x"3687", x"3689", 
    x"368c", x"368f", x"3692", x"3695", x"3698", x"369a", x"369d", x"36a0", 
    x"36a3", x"36a6", x"36a9", x"36ab", x"36ae", x"36b1", x"36b4", x"36b7", 
    x"36ba", x"36bd", x"36bf", x"36c2", x"36c5", x"36c8", x"36cb", x"36ce", 
    x"36d0", x"36d3", x"36d6", x"36d9", x"36dc", x"36df", x"36e1", x"36e4", 
    x"36e7", x"36ea", x"36ed", x"36f0", x"36f2", x"36f5", x"36f8", x"36fb", 
    x"36fe", x"3701", x"3703", x"3706", x"3709", x"370c", x"370f", x"3712", 
    x"3715", x"3717", x"371a", x"371d", x"3720", x"3723", x"3726", x"3728", 
    x"372b", x"372e", x"3731", x"3734", x"3737", x"3739", x"373c", x"373f", 
    x"3742", x"3745", x"3748", x"374a", x"374d", x"3750", x"3753", x"3756", 
    x"3759", x"375b", x"375e", x"3761", x"3764", x"3767", x"376a", x"376c", 
    x"376f", x"3772", x"3775", x"3778", x"377b", x"377d", x"3780", x"3783", 
    x"3786", x"3789", x"378b", x"378e", x"3791", x"3794", x"3797", x"379a", 
    x"379c", x"379f", x"37a2", x"37a5", x"37a8", x"37ab", x"37ad", x"37b0", 
    x"37b3", x"37b6", x"37b9", x"37bc", x"37be", x"37c1", x"37c4", x"37c7", 
    x"37ca", x"37cd", x"37cf", x"37d2", x"37d5", x"37d8", x"37db", x"37de", 
    x"37e0", x"37e3", x"37e6", x"37e9", x"37ec", x"37ee", x"37f1", x"37f4", 
    x"37f7", x"37fa", x"37fd", x"37ff", x"3802", x"3805", x"3808", x"380b", 
    x"380e", x"3810", x"3813", x"3816", x"3819", x"381c", x"381e", x"3821", 
    x"3824", x"3827", x"382a", x"382d", x"382f", x"3832", x"3835", x"3838", 
    x"383b", x"383e", x"3840", x"3843", x"3846", x"3849", x"384c", x"384e", 
    x"3851", x"3854", x"3857", x"385a", x"385d", x"385f", x"3862", x"3865", 
    x"3868", x"386b", x"386d", x"3870", x"3873", x"3876", x"3879", x"387c", 
    x"387e", x"3881", x"3884", x"3887", x"388a", x"388d", x"388f", x"3892", 
    x"3895", x"3898", x"389b", x"389d", x"38a0", x"38a3", x"38a6", x"38a9", 
    x"38ab", x"38ae", x"38b1", x"38b4", x"38b7", x"38ba", x"38bc", x"38bf", 
    x"38c2", x"38c5", x"38c8", x"38ca", x"38cd", x"38d0", x"38d3", x"38d6", 
    x"38d9", x"38db", x"38de", x"38e1", x"38e4", x"38e7", x"38e9", x"38ec", 
    x"38ef", x"38f2", x"38f5", x"38f8", x"38fa", x"38fd", x"3900", x"3903", 
    x"3906", x"3908", x"390b", x"390e", x"3911", x"3914", x"3916", x"3919", 
    x"391c", x"391f", x"3922", x"3924", x"3927", x"392a", x"392d", x"3930", 
    x"3933", x"3935", x"3938", x"393b", x"393e", x"3941", x"3943", x"3946", 
    x"3949", x"394c", x"394f", x"3951", x"3954", x"3957", x"395a", x"395d", 
    x"3960", x"3962", x"3965", x"3968", x"396b", x"396e", x"3970", x"3973", 
    x"3976", x"3979", x"397c", x"397e", x"3981", x"3984", x"3987", x"398a", 
    x"398c", x"398f", x"3992", x"3995", x"3998", x"399a", x"399d", x"39a0", 
    x"39a3", x"39a6", x"39a8", x"39ab", x"39ae", x"39b1", x"39b4", x"39b6", 
    x"39b9", x"39bc", x"39bf", x"39c2", x"39c5", x"39c7", x"39ca", x"39cd", 
    x"39d0", x"39d3", x"39d5", x"39d8", x"39db", x"39de", x"39e1", x"39e3", 
    x"39e6", x"39e9", x"39ec", x"39ef", x"39f1", x"39f4", x"39f7", x"39fa", 
    x"39fd", x"39ff", x"3a02", x"3a05", x"3a08", x"3a0b", x"3a0d", x"3a10", 
    x"3a13", x"3a16", x"3a19", x"3a1b", x"3a1e", x"3a21", x"3a24", x"3a27", 
    x"3a29", x"3a2c", x"3a2f", x"3a32", x"3a35", x"3a37", x"3a3a", x"3a3d", 
    x"3a40", x"3a43", x"3a45", x"3a48", x"3a4b", x"3a4e", x"3a51", x"3a53", 
    x"3a56", x"3a59", x"3a5c", x"3a5e", x"3a61", x"3a64", x"3a67", x"3a6a", 
    x"3a6c", x"3a6f", x"3a72", x"3a75", x"3a78", x"3a7a", x"3a7d", x"3a80", 
    x"3a83", x"3a86", x"3a88", x"3a8b", x"3a8e", x"3a91", x"3a94", x"3a96", 
    x"3a99", x"3a9c", x"3a9f", x"3aa2", x"3aa4", x"3aa7", x"3aaa", x"3aad", 
    x"3ab0", x"3ab2", x"3ab5", x"3ab8", x"3abb", x"3abd", x"3ac0", x"3ac3", 
    x"3ac6", x"3ac9", x"3acb", x"3ace", x"3ad1", x"3ad4", x"3ad7", x"3ad9", 
    x"3adc", x"3adf", x"3ae2", x"3ae5", x"3ae7", x"3aea", x"3aed", x"3af0", 
    x"3af2", x"3af5", x"3af8", x"3afb", x"3afe", x"3b00", x"3b03", x"3b06", 
    x"3b09", x"3b0c", x"3b0e", x"3b11", x"3b14", x"3b17", x"3b19", x"3b1c", 
    x"3b1f", x"3b22", x"3b25", x"3b27", x"3b2a", x"3b2d", x"3b30", x"3b33", 
    x"3b35", x"3b38", x"3b3b", x"3b3e", x"3b40", x"3b43", x"3b46", x"3b49", 
    x"3b4c", x"3b4e", x"3b51", x"3b54", x"3b57", x"3b5a", x"3b5c", x"3b5f", 
    x"3b62", x"3b65", x"3b67", x"3b6a", x"3b6d", x"3b70", x"3b73", x"3b75", 
    x"3b78", x"3b7b", x"3b7e", x"3b81", x"3b83", x"3b86", x"3b89", x"3b8c", 
    x"3b8e", x"3b91", x"3b94", x"3b97", x"3b9a", x"3b9c", x"3b9f", x"3ba2", 
    x"3ba5", x"3ba7", x"3baa", x"3bad", x"3bb0", x"3bb3", x"3bb5", x"3bb8", 
    x"3bbb", x"3bbe", x"3bc0", x"3bc3", x"3bc6", x"3bc9", x"3bcc", x"3bce", 
    x"3bd1", x"3bd4", x"3bd7", x"3bd9", x"3bdc", x"3bdf", x"3be2", x"3be5", 
    x"3be7", x"3bea", x"3bed", x"3bf0", x"3bf2", x"3bf5", x"3bf8", x"3bfb", 
    x"3bfe", x"3c00", x"3c03", x"3c06", x"3c09", x"3c0b", x"3c0e", x"3c11", 
    x"3c14", x"3c16", x"3c19", x"3c1c", x"3c1f", x"3c22", x"3c24", x"3c27", 
    x"3c2a", x"3c2d", x"3c2f", x"3c32", x"3c35", x"3c38", x"3c3b", x"3c3d", 
    x"3c40", x"3c43", x"3c46", x"3c48", x"3c4b", x"3c4e", x"3c51", x"3c53", 
    x"3c56", x"3c59", x"3c5c", x"3c5f", x"3c61", x"3c64", x"3c67", x"3c6a", 
    x"3c6c", x"3c6f", x"3c72", x"3c75", x"3c77", x"3c7a", x"3c7d", x"3c80", 
    x"3c83", x"3c85", x"3c88", x"3c8b", x"3c8e", x"3c90", x"3c93", x"3c96", 
    x"3c99", x"3c9b", x"3c9e", x"3ca1", x"3ca4", x"3ca7", x"3ca9", x"3cac", 
    x"3caf", x"3cb2", x"3cb4", x"3cb7", x"3cba", x"3cbd", x"3cbf", x"3cc2", 
    x"3cc5", x"3cc8", x"3cca", x"3ccd", x"3cd0", x"3cd3", x"3cd6", x"3cd8", 
    x"3cdb", x"3cde", x"3ce1", x"3ce3", x"3ce6", x"3ce9", x"3cec", x"3cee", 
    x"3cf1", x"3cf4", x"3cf7", x"3cf9", x"3cfc", x"3cff", x"3d02", x"3d05", 
    x"3d07", x"3d0a", x"3d0d", x"3d10", x"3d12", x"3d15", x"3d18", x"3d1b", 
    x"3d1d", x"3d20", x"3d23", x"3d26", x"3d28", x"3d2b", x"3d2e", x"3d31", 
    x"3d33", x"3d36", x"3d39", x"3d3c", x"3d3e", x"3d41", x"3d44", x"3d47", 
    x"3d4a", x"3d4c", x"3d4f", x"3d52", x"3d55", x"3d57", x"3d5a", x"3d5d", 
    x"3d60", x"3d62", x"3d65", x"3d68", x"3d6b", x"3d6d", x"3d70", x"3d73", 
    x"3d76", x"3d78", x"3d7b", x"3d7e", x"3d81", x"3d83", x"3d86", x"3d89", 
    x"3d8c", x"3d8e", x"3d91", x"3d94", x"3d97", x"3d99", x"3d9c", x"3d9f", 
    x"3da2", x"3da4", x"3da7", x"3daa", x"3dad", x"3daf", x"3db2", x"3db5", 
    x"3db8", x"3dba", x"3dbd", x"3dc0", x"3dc3", x"3dc5", x"3dc8", x"3dcb", 
    x"3dce", x"3dd0", x"3dd3", x"3dd6", x"3dd9", x"3ddb", x"3dde", x"3de1", 
    x"3de4", x"3de6", x"3de9", x"3dec", x"3def", x"3df1", x"3df4", x"3df7", 
    x"3dfa", x"3dfc", x"3dff", x"3e02", x"3e05", x"3e07", x"3e0a", x"3e0d", 
    x"3e10", x"3e12", x"3e15", x"3e18", x"3e1b", x"3e1d", x"3e20", x"3e23", 
    x"3e26", x"3e28", x"3e2b", x"3e2e", x"3e31", x"3e33", x"3e36", x"3e39", 
    x"3e3c", x"3e3e", x"3e41", x"3e44", x"3e47", x"3e49", x"3e4c", x"3e4f", 
    x"3e52", x"3e54", x"3e57", x"3e5a", x"3e5d", x"3e5f", x"3e62", x"3e65", 
    x"3e68", x"3e6a", x"3e6d", x"3e70", x"3e73", x"3e75", x"3e78", x"3e7b", 
    x"3e7d", x"3e80", x"3e83", x"3e86", x"3e88", x"3e8b", x"3e8e", x"3e91", 
    x"3e93", x"3e96", x"3e99", x"3e9c", x"3e9e", x"3ea1", x"3ea4", x"3ea7", 
    x"3ea9", x"3eac", x"3eaf", x"3eb2", x"3eb4", x"3eb7", x"3eba", x"3ebd", 
    x"3ebf", x"3ec2", x"3ec5", x"3ec7", x"3eca", x"3ecd", x"3ed0", x"3ed2", 
    x"3ed5", x"3ed8", x"3edb", x"3edd", x"3ee0", x"3ee3", x"3ee6", x"3ee8", 
    x"3eeb", x"3eee", x"3ef1", x"3ef3", x"3ef6", x"3ef9", x"3efb", x"3efe", 
    x"3f01", x"3f04", x"3f06", x"3f09", x"3f0c", x"3f0f", x"3f11", x"3f14", 
    x"3f17", x"3f1a", x"3f1c", x"3f1f", x"3f22", x"3f24", x"3f27", x"3f2a", 
    x"3f2d", x"3f2f", x"3f32", x"3f35", x"3f38", x"3f3a", x"3f3d", x"3f40", 
    x"3f43", x"3f45", x"3f48", x"3f4b", x"3f4d", x"3f50", x"3f53", x"3f56", 
    x"3f58", x"3f5b", x"3f5e", x"3f61", x"3f63", x"3f66", x"3f69", x"3f6b", 
    x"3f6e", x"3f71", x"3f74", x"3f76", x"3f79", x"3f7c", x"3f7f", x"3f81", 
    x"3f84", x"3f87", x"3f89", x"3f8c", x"3f8f", x"3f92", x"3f94", x"3f97", 
    x"3f9a", x"3f9d", x"3f9f", x"3fa2", x"3fa5", x"3fa7", x"3faa", x"3fad", 
    x"3fb0", x"3fb2", x"3fb5", x"3fb8", x"3fbb", x"3fbd", x"3fc0", x"3fc3", 
    x"3fc5", x"3fc8", x"3fcb", x"3fce", x"3fd0", x"3fd3", x"3fd6", x"3fd8", 
    x"3fdb", x"3fde", x"3fe1", x"3fe3", x"3fe6", x"3fe9", x"3fec", x"3fee", 
    x"3ff1", x"3ff4", x"3ff6", x"3ff9", x"3ffc", x"3fff", x"4001", x"4004", 
    x"4007", x"4009", x"400c", x"400f", x"4012", x"4014", x"4017", x"401a", 
    x"401d", x"401f", x"4022", x"4025", x"4027", x"402a", x"402d", x"4030", 
    x"4032", x"4035", x"4038", x"403a", x"403d", x"4040", x"4043", x"4045", 
    x"4048", x"404b", x"404d", x"4050", x"4053", x"4056", x"4058", x"405b", 
    x"405e", x"4060", x"4063", x"4066", x"4069", x"406b", x"406e", x"4071", 
    x"4073", x"4076", x"4079", x"407c", x"407e", x"4081", x"4084", x"4086", 
    x"4089", x"408c", x"408f", x"4091", x"4094", x"4097", x"4099", x"409c", 
    x"409f", x"40a2", x"40a4", x"40a7", x"40aa", x"40ac", x"40af", x"40b2", 
    x"40b5", x"40b7", x"40ba", x"40bd", x"40bf", x"40c2", x"40c5", x"40c8", 
    x"40ca", x"40cd", x"40d0", x"40d2", x"40d5", x"40d8", x"40da", x"40dd", 
    x"40e0", x"40e3", x"40e5", x"40e8", x"40eb", x"40ed", x"40f0", x"40f3", 
    x"40f6", x"40f8", x"40fb", x"40fe", x"4100", x"4103", x"4106", x"4108", 
    x"410b", x"410e", x"4111", x"4113", x"4116", x"4119", x"411b", x"411e", 
    x"4121", x"4124", x"4126", x"4129", x"412c", x"412e", x"4131", x"4134", 
    x"4136", x"4139", x"413c", x"413f", x"4141", x"4144", x"4147", x"4149", 
    x"414c", x"414f", x"4151", x"4154", x"4157", x"415a", x"415c", x"415f", 
    x"4162", x"4164", x"4167", x"416a", x"416d", x"416f", x"4172", x"4175", 
    x"4177", x"417a", x"417d", x"417f", x"4182", x"4185", x"4187", x"418a", 
    x"418d", x"4190", x"4192", x"4195", x"4198", x"419a", x"419d", x"41a0", 
    x"41a2", x"41a5", x"41a8", x"41ab", x"41ad", x"41b0", x"41b3", x"41b5", 
    x"41b8", x"41bb", x"41bd", x"41c0", x"41c3", x"41c6", x"41c8", x"41cb", 
    x"41ce", x"41d0", x"41d3", x"41d6", x"41d8", x"41db", x"41de", x"41e0", 
    x"41e3", x"41e6", x"41e9", x"41eb", x"41ee", x"41f1", x"41f3", x"41f6", 
    x"41f9", x"41fb", x"41fe", x"4201", x"4203", x"4206", x"4209", x"420c", 
    x"420e", x"4211", x"4214", x"4216", x"4219", x"421c", x"421e", x"4221", 
    x"4224", x"4226", x"4229", x"422c", x"422f", x"4231", x"4234", x"4237", 
    x"4239", x"423c", x"423f", x"4241", x"4244", x"4247", x"4249", x"424c", 
    x"424f", x"4251", x"4254", x"4257", x"425a", x"425c", x"425f", x"4262", 
    x"4264", x"4267", x"426a", x"426c", x"426f", x"4272", x"4274", x"4277", 
    x"427a", x"427c", x"427f", x"4282", x"4284", x"4287", x"428a", x"428d", 
    x"428f", x"4292", x"4295", x"4297", x"429a", x"429d", x"429f", x"42a2", 
    x"42a5", x"42a7", x"42aa", x"42ad", x"42af", x"42b2", x"42b5", x"42b7", 
    x"42ba", x"42bd", x"42bf", x"42c2", x"42c5", x"42c8", x"42ca", x"42cd", 
    x"42d0", x"42d2", x"42d5", x"42d8", x"42da", x"42dd", x"42e0", x"42e2", 
    x"42e5", x"42e8", x"42ea", x"42ed", x"42f0", x"42f2", x"42f5", x"42f8", 
    x"42fa", x"42fd", x"4300", x"4302", x"4305", x"4308", x"430a", x"430d", 
    x"4310", x"4313", x"4315", x"4318", x"431b", x"431d", x"4320", x"4323", 
    x"4325", x"4328", x"432b", x"432d", x"4330", x"4333", x"4335", x"4338", 
    x"433b", x"433d", x"4340", x"4343", x"4345", x"4348", x"434b", x"434d", 
    x"4350", x"4353", x"4355", x"4358", x"435b", x"435d", x"4360", x"4363", 
    x"4365", x"4368", x"436b", x"436d", x"4370", x"4373", x"4375", x"4378", 
    x"437b", x"437d", x"4380", x"4383", x"4385", x"4388", x"438b", x"438d", 
    x"4390", x"4393", x"4395", x"4398", x"439b", x"439d", x"43a0", x"43a3", 
    x"43a5", x"43a8", x"43ab", x"43ad", x"43b0", x"43b3", x"43b5", x"43b8", 
    x"43bb", x"43bd", x"43c0", x"43c3", x"43c5", x"43c8", x"43cb", x"43cd", 
    x"43d0", x"43d3", x"43d5", x"43d8", x"43db", x"43dd", x"43e0", x"43e3", 
    x"43e5", x"43e8", x"43eb", x"43ed", x"43f0", x"43f3", x"43f5", x"43f8", 
    x"43fb", x"43fd", x"4400", x"4403", x"4405", x"4408", x"440b", x"440d", 
    x"4410", x"4413", x"4415", x"4418", x"441b", x"441d", x"4420", x"4423", 
    x"4425", x"4428", x"442b", x"442d", x"4430", x"4433", x"4435", x"4438", 
    x"443b", x"443d", x"4440", x"4442", x"4445", x"4448", x"444a", x"444d", 
    x"4450", x"4452", x"4455", x"4458", x"445a", x"445d", x"4460", x"4462", 
    x"4465", x"4468", x"446a", x"446d", x"4470", x"4472", x"4475", x"4478", 
    x"447a", x"447d", x"4480", x"4482", x"4485", x"4488", x"448a", x"448d", 
    x"448f", x"4492", x"4495", x"4497", x"449a", x"449d", x"449f", x"44a2", 
    x"44a5", x"44a7", x"44aa", x"44ad", x"44af", x"44b2", x"44b5", x"44b7", 
    x"44ba", x"44bd", x"44bf", x"44c2", x"44c5", x"44c7", x"44ca", x"44cc", 
    x"44cf", x"44d2", x"44d4", x"44d7", x"44da", x"44dc", x"44df", x"44e2", 
    x"44e4", x"44e7", x"44ea", x"44ec", x"44ef", x"44f2", x"44f4", x"44f7", 
    x"44f9", x"44fc", x"44ff", x"4501", x"4504", x"4507", x"4509", x"450c", 
    x"450f", x"4511", x"4514", x"4517", x"4519", x"451c", x"451f", x"4521", 
    x"4524", x"4526", x"4529", x"452c", x"452e", x"4531", x"4534", x"4536", 
    x"4539", x"453c", x"453e", x"4541", x"4544", x"4546", x"4549", x"454b", 
    x"454e", x"4551", x"4553", x"4556", x"4559", x"455b", x"455e", x"4561", 
    x"4563", x"4566", x"4568", x"456b", x"456e", x"4570", x"4573", x"4576", 
    x"4578", x"457b", x"457e", x"4580", x"4583", x"4586", x"4588", x"458b", 
    x"458d", x"4590", x"4593", x"4595", x"4598", x"459b", x"459d", x"45a0", 
    x"45a3", x"45a5", x"45a8", x"45aa", x"45ad", x"45b0", x"45b2", x"45b5", 
    x"45b8", x"45ba", x"45bd", x"45bf", x"45c2", x"45c5", x"45c7", x"45ca", 
    x"45cd", x"45cf", x"45d2", x"45d5", x"45d7", x"45da", x"45dc", x"45df", 
    x"45e2", x"45e4", x"45e7", x"45ea", x"45ec", x"45ef", x"45f2", x"45f4", 
    x"45f7", x"45f9", x"45fc", x"45ff", x"4601", x"4604", x"4607", x"4609", 
    x"460c", x"460e", x"4611", x"4614", x"4616", x"4619", x"461c", x"461e", 
    x"4621", x"4623", x"4626", x"4629", x"462b", x"462e", x"4631", x"4633", 
    x"4636", x"4638", x"463b", x"463e", x"4640", x"4643", x"4646", x"4648", 
    x"464b", x"464d", x"4650", x"4653", x"4655", x"4658", x"465b", x"465d", 
    x"4660", x"4662", x"4665", x"4668", x"466a", x"466d", x"4670", x"4672", 
    x"4675", x"4677", x"467a", x"467d", x"467f", x"4682", x"4685", x"4687", 
    x"468a", x"468c", x"468f", x"4692", x"4694", x"4697", x"469a", x"469c", 
    x"469f", x"46a1", x"46a4", x"46a7", x"46a9", x"46ac", x"46af", x"46b1", 
    x"46b4", x"46b6", x"46b9", x"46bc", x"46be", x"46c1", x"46c3", x"46c6", 
    x"46c9", x"46cb", x"46ce", x"46d1", x"46d3", x"46d6", x"46d8", x"46db", 
    x"46de", x"46e0", x"46e3", x"46e5", x"46e8", x"46eb", x"46ed", x"46f0", 
    x"46f3", x"46f5", x"46f8", x"46fa", x"46fd", x"4700", x"4702", x"4705", 
    x"4707", x"470a", x"470d", x"470f", x"4712", x"4715", x"4717", x"471a", 
    x"471c", x"471f", x"4722", x"4724", x"4727", x"4729", x"472c", x"472f", 
    x"4731", x"4734", x"4736", x"4739", x"473c", x"473e", x"4741", x"4744", 
    x"4746", x"4749", x"474b", x"474e", x"4751", x"4753", x"4756", x"4758", 
    x"475b", x"475e", x"4760", x"4763", x"4765", x"4768", x"476b", x"476d", 
    x"4770", x"4772", x"4775", x"4778", x"477a", x"477d", x"4780", x"4782", 
    x"4785", x"4787", x"478a", x"478d", x"478f", x"4792", x"4794", x"4797", 
    x"479a", x"479c", x"479f", x"47a1", x"47a4", x"47a7", x"47a9", x"47ac", 
    x"47ae", x"47b1", x"47b4", x"47b6", x"47b9", x"47bb", x"47be", x"47c1", 
    x"47c3", x"47c6", x"47c8", x"47cb", x"47ce", x"47d0", x"47d3", x"47d5", 
    x"47d8", x"47db", x"47dd", x"47e0", x"47e2", x"47e5", x"47e8", x"47ea", 
    x"47ed", x"47ef", x"47f2", x"47f5", x"47f7", x"47fa", x"47fc", x"47ff", 
    x"4802", x"4804", x"4807", x"4809", x"480c", x"480f", x"4811", x"4814", 
    x"4816", x"4819", x"481c", x"481e", x"4821", x"4823", x"4826", x"4829", 
    x"482b", x"482e", x"4830", x"4833", x"4835", x"4838", x"483b", x"483d", 
    x"4840", x"4842", x"4845", x"4848", x"484a", x"484d", x"484f", x"4852", 
    x"4855", x"4857", x"485a", x"485c", x"485f", x"4862", x"4864", x"4867", 
    x"4869", x"486c", x"486f", x"4871", x"4874", x"4876", x"4879", x"487b", 
    x"487e", x"4881", x"4883", x"4886", x"4888", x"488b", x"488e", x"4890", 
    x"4893", x"4895", x"4898", x"489b", x"489d", x"48a0", x"48a2", x"48a5", 
    x"48a7", x"48aa", x"48ad", x"48af", x"48b2", x"48b4", x"48b7", x"48ba", 
    x"48bc", x"48bf", x"48c1", x"48c4", x"48c6", x"48c9", x"48cc", x"48ce", 
    x"48d1", x"48d3", x"48d6", x"48d9", x"48db", x"48de", x"48e0", x"48e3", 
    x"48e5", x"48e8", x"48eb", x"48ed", x"48f0", x"48f2", x"48f5", x"48f8", 
    x"48fa", x"48fd", x"48ff", x"4902", x"4904", x"4907", x"490a", x"490c", 
    x"490f", x"4911", x"4914", x"4917", x"4919", x"491c", x"491e", x"4921", 
    x"4923", x"4926", x"4929", x"492b", x"492e", x"4930", x"4933", x"4935", 
    x"4938", x"493b", x"493d", x"4940", x"4942", x"4945", x"4947", x"494a", 
    x"494d", x"494f", x"4952", x"4954", x"4957", x"495a", x"495c", x"495f", 
    x"4961", x"4964", x"4966", x"4969", x"496c", x"496e", x"4971", x"4973", 
    x"4976", x"4978", x"497b", x"497e", x"4980", x"4983", x"4985", x"4988", 
    x"498a", x"498d", x"4990", x"4992", x"4995", x"4997", x"499a", x"499c", 
    x"499f", x"49a2", x"49a4", x"49a7", x"49a9", x"49ac", x"49ae", x"49b1", 
    x"49b4", x"49b6", x"49b9", x"49bb", x"49be", x"49c0", x"49c3", x"49c5", 
    x"49c8", x"49cb", x"49cd", x"49d0", x"49d2", x"49d5", x"49d7", x"49da", 
    x"49dd", x"49df", x"49e2", x"49e4", x"49e7", x"49e9", x"49ec", x"49ef", 
    x"49f1", x"49f4", x"49f6", x"49f9", x"49fb", x"49fe", x"4a00", x"4a03", 
    x"4a06", x"4a08", x"4a0b", x"4a0d", x"4a10", x"4a12", x"4a15", x"4a18", 
    x"4a1a", x"4a1d", x"4a1f", x"4a22", x"4a24", x"4a27", x"4a29", x"4a2c", 
    x"4a2f", x"4a31", x"4a34", x"4a36", x"4a39", x"4a3b", x"4a3e", x"4a41", 
    x"4a43", x"4a46", x"4a48", x"4a4b", x"4a4d", x"4a50", x"4a52", x"4a55", 
    x"4a58", x"4a5a", x"4a5d", x"4a5f", x"4a62", x"4a64", x"4a67", x"4a69", 
    x"4a6c", x"4a6f", x"4a71", x"4a74", x"4a76", x"4a79", x"4a7b", x"4a7e", 
    x"4a80", x"4a83", x"4a86", x"4a88", x"4a8b", x"4a8d", x"4a90", x"4a92", 
    x"4a95", x"4a97", x"4a9a", x"4a9d", x"4a9f", x"4aa2", x"4aa4", x"4aa7", 
    x"4aa9", x"4aac", x"4aae", x"4ab1", x"4ab3", x"4ab6", x"4ab9", x"4abb", 
    x"4abe", x"4ac0", x"4ac3", x"4ac5", x"4ac8", x"4aca", x"4acd", x"4ad0", 
    x"4ad2", x"4ad5", x"4ad7", x"4ada", x"4adc", x"4adf", x"4ae1", x"4ae4", 
    x"4ae6", x"4ae9", x"4aec", x"4aee", x"4af1", x"4af3", x"4af6", x"4af8", 
    x"4afb", x"4afd", x"4b00", x"4b02", x"4b05", x"4b08", x"4b0a", x"4b0d", 
    x"4b0f", x"4b12", x"4b14", x"4b17", x"4b19", x"4b1c", x"4b1e", x"4b21", 
    x"4b24", x"4b26", x"4b29", x"4b2b", x"4b2e", x"4b30", x"4b33", x"4b35", 
    x"4b38", x"4b3a", x"4b3d", x"4b40", x"4b42", x"4b45", x"4b47", x"4b4a", 
    x"4b4c", x"4b4f", x"4b51", x"4b54", x"4b56", x"4b59", x"4b5b", x"4b5e", 
    x"4b61", x"4b63", x"4b66", x"4b68", x"4b6b", x"4b6d", x"4b70", x"4b72", 
    x"4b75", x"4b77", x"4b7a", x"4b7c", x"4b7f", x"4b82", x"4b84", x"4b87", 
    x"4b89", x"4b8c", x"4b8e", x"4b91", x"4b93", x"4b96", x"4b98", x"4b9b", 
    x"4b9d", x"4ba0", x"4ba2", x"4ba5", x"4ba8", x"4baa", x"4bad", x"4baf", 
    x"4bb2", x"4bb4", x"4bb7", x"4bb9", x"4bbc", x"4bbe", x"4bc1", x"4bc3", 
    x"4bc6", x"4bc8", x"4bcb", x"4bce", x"4bd0", x"4bd3", x"4bd5", x"4bd8", 
    x"4bda", x"4bdd", x"4bdf", x"4be2", x"4be4", x"4be7", x"4be9", x"4bec", 
    x"4bee", x"4bf1", x"4bf4", x"4bf6", x"4bf9", x"4bfb", x"4bfe", x"4c00", 
    x"4c03", x"4c05", x"4c08", x"4c0a", x"4c0d", x"4c0f", x"4c12", x"4c14", 
    x"4c17", x"4c19", x"4c1c", x"4c1e", x"4c21", x"4c24", x"4c26", x"4c29", 
    x"4c2b", x"4c2e", x"4c30", x"4c33", x"4c35", x"4c38", x"4c3a", x"4c3d", 
    x"4c3f", x"4c42", x"4c44", x"4c47", x"4c49", x"4c4c", x"4c4e", x"4c51", 
    x"4c53", x"4c56", x"4c59", x"4c5b", x"4c5e", x"4c60", x"4c63", x"4c65", 
    x"4c68", x"4c6a", x"4c6d", x"4c6f", x"4c72", x"4c74", x"4c77", x"4c79", 
    x"4c7c", x"4c7e", x"4c81", x"4c83", x"4c86", x"4c88", x"4c8b", x"4c8d", 
    x"4c90", x"4c92", x"4c95", x"4c97", x"4c9a", x"4c9d", x"4c9f", x"4ca2", 
    x"4ca4", x"4ca7", x"4ca9", x"4cac", x"4cae", x"4cb1", x"4cb3", x"4cb6", 
    x"4cb8", x"4cbb", x"4cbd", x"4cc0", x"4cc2", x"4cc5", x"4cc7", x"4cca", 
    x"4ccc", x"4ccf", x"4cd1", x"4cd4", x"4cd6", x"4cd9", x"4cdb", x"4cde", 
    x"4ce0", x"4ce3", x"4ce5", x"4ce8", x"4cea", x"4ced", x"4cef", x"4cf2", 
    x"4cf4", x"4cf7", x"4cfa", x"4cfc", x"4cff", x"4d01", x"4d04", x"4d06", 
    x"4d09", x"4d0b", x"4d0e", x"4d10", x"4d13", x"4d15", x"4d18", x"4d1a", 
    x"4d1d", x"4d1f", x"4d22", x"4d24", x"4d27", x"4d29", x"4d2c", x"4d2e", 
    x"4d31", x"4d33", x"4d36", x"4d38", x"4d3b", x"4d3d", x"4d40", x"4d42", 
    x"4d45", x"4d47", x"4d4a", x"4d4c", x"4d4f", x"4d51", x"4d54", x"4d56", 
    x"4d59", x"4d5b", x"4d5e", x"4d60", x"4d63", x"4d65", x"4d68", x"4d6a", 
    x"4d6d", x"4d6f", x"4d72", x"4d74", x"4d77", x"4d79", x"4d7c", x"4d7e", 
    x"4d81", x"4d83", x"4d86", x"4d88", x"4d8b", x"4d8d", x"4d90", x"4d92", 
    x"4d95", x"4d97", x"4d9a", x"4d9c", x"4d9f", x"4da1", x"4da4", x"4da6", 
    x"4da9", x"4dab", x"4dae", x"4db0", x"4db3", x"4db5", x"4db8", x"4dba", 
    x"4dbd", x"4dbf", x"4dc2", x"4dc4", x"4dc7", x"4dc9", x"4dcc", x"4dce", 
    x"4dd1", x"4dd3", x"4dd6", x"4dd8", x"4ddb", x"4ddd", x"4de0", x"4de2", 
    x"4de5", x"4de7", x"4dea", x"4dec", x"4def", x"4df1", x"4df4", x"4df6", 
    x"4df9", x"4dfb", x"4dfe", x"4e00", x"4e03", x"4e05", x"4e08", x"4e0a", 
    x"4e0d", x"4e0f", x"4e11", x"4e14", x"4e16", x"4e19", x"4e1b", x"4e1e", 
    x"4e20", x"4e23", x"4e25", x"4e28", x"4e2a", x"4e2d", x"4e2f", x"4e32", 
    x"4e34", x"4e37", x"4e39", x"4e3c", x"4e3e", x"4e41", x"4e43", x"4e46", 
    x"4e48", x"4e4b", x"4e4d", x"4e50", x"4e52", x"4e55", x"4e57", x"4e5a", 
    x"4e5c", x"4e5f", x"4e61", x"4e64", x"4e66", x"4e68", x"4e6b", x"4e6d", 
    x"4e70", x"4e72", x"4e75", x"4e77", x"4e7a", x"4e7c", x"4e7f", x"4e81", 
    x"4e84", x"4e86", x"4e89", x"4e8b", x"4e8e", x"4e90", x"4e93", x"4e95", 
    x"4e98", x"4e9a", x"4e9d", x"4e9f", x"4ea2", x"4ea4", x"4ea7", x"4ea9", 
    x"4eab", x"4eae", x"4eb0", x"4eb3", x"4eb5", x"4eb8", x"4eba", x"4ebd", 
    x"4ebf", x"4ec2", x"4ec4", x"4ec7", x"4ec9", x"4ecc", x"4ece", x"4ed1", 
    x"4ed3", x"4ed6", x"4ed8", x"4edb", x"4edd", x"4edf", x"4ee2", x"4ee4", 
    x"4ee7", x"4ee9", x"4eec", x"4eee", x"4ef1", x"4ef3", x"4ef6", x"4ef8", 
    x"4efb", x"4efd", x"4f00", x"4f02", x"4f05", x"4f07", x"4f0a", x"4f0c", 
    x"4f0e", x"4f11", x"4f13", x"4f16", x"4f18", x"4f1b", x"4f1d", x"4f20", 
    x"4f22", x"4f25", x"4f27", x"4f2a", x"4f2c", x"4f2f", x"4f31", x"4f33", 
    x"4f36", x"4f38", x"4f3b", x"4f3d", x"4f40", x"4f42", x"4f45", x"4f47", 
    x"4f4a", x"4f4c", x"4f4f", x"4f51", x"4f54", x"4f56", x"4f58", x"4f5b", 
    x"4f5d", x"4f60", x"4f62", x"4f65", x"4f67", x"4f6a", x"4f6c", x"4f6f", 
    x"4f71", x"4f74", x"4f76", x"4f79", x"4f7b", x"4f7d", x"4f80", x"4f82", 
    x"4f85", x"4f87", x"4f8a", x"4f8c", x"4f8f", x"4f91", x"4f94", x"4f96", 
    x"4f99", x"4f9b", x"4f9d", x"4fa0", x"4fa2", x"4fa5", x"4fa7", x"4faa", 
    x"4fac", x"4faf", x"4fb1", x"4fb4", x"4fb6", x"4fb8", x"4fbb", x"4fbd", 
    x"4fc0", x"4fc2", x"4fc5", x"4fc7", x"4fca", x"4fcc", x"4fcf", x"4fd1", 
    x"4fd4", x"4fd6", x"4fd8", x"4fdb", x"4fdd", x"4fe0", x"4fe2", x"4fe5", 
    x"4fe7", x"4fea", x"4fec", x"4fef", x"4ff1", x"4ff3", x"4ff6", x"4ff8", 
    x"4ffb", x"4ffd", x"5000", x"5002", x"5005", x"5007", x"5009", x"500c", 
    x"500e", x"5011", x"5013", x"5016", x"5018", x"501b", x"501d", x"5020", 
    x"5022", x"5024", x"5027", x"5029", x"502c", x"502e", x"5031", x"5033", 
    x"5036", x"5038", x"503a", x"503d", x"503f", x"5042", x"5044", x"5047", 
    x"5049", x"504c", x"504e", x"5050", x"5053", x"5055", x"5058", x"505a", 
    x"505d", x"505f", x"5062", x"5064", x"5067", x"5069", x"506b", x"506e", 
    x"5070", x"5073", x"5075", x"5078", x"507a", x"507c", x"507f", x"5081", 
    x"5084", x"5086", x"5089", x"508b", x"508e", x"5090", x"5092", x"5095", 
    x"5097", x"509a", x"509c", x"509f", x"50a1", x"50a4", x"50a6", x"50a8", 
    x"50ab", x"50ad", x"50b0", x"50b2", x"50b5", x"50b7", x"50ba", x"50bc", 
    x"50be", x"50c1", x"50c3", x"50c6", x"50c8", x"50cb", x"50cd", x"50cf", 
    x"50d2", x"50d4", x"50d7", x"50d9", x"50dc", x"50de", x"50e0", x"50e3", 
    x"50e5", x"50e8", x"50ea", x"50ed", x"50ef", x"50f2", x"50f4", x"50f6", 
    x"50f9", x"50fb", x"50fe", x"5100", x"5103", x"5105", x"5107", x"510a", 
    x"510c", x"510f", x"5111", x"5114", x"5116", x"5118", x"511b", x"511d", 
    x"5120", x"5122", x"5125", x"5127", x"5129", x"512c", x"512e", x"5131", 
    x"5133", x"5136", x"5138", x"513a", x"513d", x"513f", x"5142", x"5144", 
    x"5147", x"5149", x"514b", x"514e", x"5150", x"5153", x"5155", x"5158", 
    x"515a", x"515c", x"515f", x"5161", x"5164", x"5166", x"5169", x"516b", 
    x"516d", x"5170", x"5172", x"5175", x"5177", x"517a", x"517c", x"517e", 
    x"5181", x"5183", x"5186", x"5188", x"518a", x"518d", x"518f", x"5192", 
    x"5194", x"5197", x"5199", x"519b", x"519e", x"51a0", x"51a3", x"51a5", 
    x"51a8", x"51aa", x"51ac", x"51af", x"51b1", x"51b4", x"51b6", x"51b8", 
    x"51bb", x"51bd", x"51c0", x"51c2", x"51c5", x"51c7", x"51c9", x"51cc", 
    x"51ce", x"51d1", x"51d3", x"51d5", x"51d8", x"51da", x"51dd", x"51df", 
    x"51e2", x"51e4", x"51e6", x"51e9", x"51eb", x"51ee", x"51f0", x"51f2", 
    x"51f5", x"51f7", x"51fa", x"51fc", x"51fe", x"5201", x"5203", x"5206", 
    x"5208", x"520b", x"520d", x"520f", x"5212", x"5214", x"5217", x"5219", 
    x"521b", x"521e", x"5220", x"5223", x"5225", x"5227", x"522a", x"522c", 
    x"522f", x"5231", x"5233", x"5236", x"5238", x"523b", x"523d", x"5240", 
    x"5242", x"5244", x"5247", x"5249", x"524c", x"524e", x"5250", x"5253", 
    x"5255", x"5258", x"525a", x"525c", x"525f", x"5261", x"5264", x"5266", 
    x"5268", x"526b", x"526d", x"5270", x"5272", x"5274", x"5277", x"5279", 
    x"527c", x"527e", x"5280", x"5283", x"5285", x"5288", x"528a", x"528c", 
    x"528f", x"5291", x"5294", x"5296", x"5298", x"529b", x"529d", x"52a0", 
    x"52a2", x"52a4", x"52a7", x"52a9", x"52ac", x"52ae", x"52b0", x"52b3", 
    x"52b5", x"52b8", x"52ba", x"52bc", x"52bf", x"52c1", x"52c4", x"52c6", 
    x"52c8", x"52cb", x"52cd", x"52d0", x"52d2", x"52d4", x"52d7", x"52d9", 
    x"52dc", x"52de", x"52e0", x"52e3", x"52e5", x"52e8", x"52ea", x"52ec", 
    x"52ef", x"52f1", x"52f4", x"52f6", x"52f8", x"52fb", x"52fd", x"52ff", 
    x"5302", x"5304", x"5307", x"5309", x"530b", x"530e", x"5310", x"5313", 
    x"5315", x"5317", x"531a", x"531c", x"531f", x"5321", x"5323", x"5326", 
    x"5328", x"532a", x"532d", x"532f", x"5332", x"5334", x"5336", x"5339", 
    x"533b", x"533e", x"5340", x"5342", x"5345", x"5347", x"534a", x"534c", 
    x"534e", x"5351", x"5353", x"5355", x"5358", x"535a", x"535d", x"535f", 
    x"5361", x"5364", x"5366", x"5369", x"536b", x"536d", x"5370", x"5372", 
    x"5374", x"5377", x"5379", x"537c", x"537e", x"5380", x"5383", x"5385", 
    x"5387", x"538a", x"538c", x"538f", x"5391", x"5393", x"5396", x"5398", 
    x"539b", x"539d", x"539f", x"53a2", x"53a4", x"53a6", x"53a9", x"53ab", 
    x"53ae", x"53b0", x"53b2", x"53b5", x"53b7", x"53b9", x"53bc", x"53be", 
    x"53c1", x"53c3", x"53c5", x"53c8", x"53ca", x"53cc", x"53cf", x"53d1", 
    x"53d4", x"53d6", x"53d8", x"53db", x"53dd", x"53df", x"53e2", x"53e4", 
    x"53e7", x"53e9", x"53eb", x"53ee", x"53f0", x"53f2", x"53f5", x"53f7", 
    x"53fa", x"53fc", x"53fe", x"5401", x"5403", x"5405", x"5408", x"540a", 
    x"540c", x"540f", x"5411", x"5414", x"5416", x"5418", x"541b", x"541d", 
    x"541f", x"5422", x"5424", x"5427", x"5429", x"542b", x"542e", x"5430", 
    x"5432", x"5435", x"5437", x"5439", x"543c", x"543e", x"5441", x"5443", 
    x"5445", x"5448", x"544a", x"544c", x"544f", x"5451", x"5453", x"5456", 
    x"5458", x"545b", x"545d", x"545f", x"5462", x"5464", x"5466", x"5469", 
    x"546b", x"546d", x"5470", x"5472", x"5475", x"5477", x"5479", x"547c", 
    x"547e", x"5480", x"5483", x"5485", x"5487", x"548a", x"548c", x"548e", 
    x"5491", x"5493", x"5496", x"5498", x"549a", x"549d", x"549f", x"54a1", 
    x"54a4", x"54a6", x"54a8", x"54ab", x"54ad", x"54af", x"54b2", x"54b4", 
    x"54b7", x"54b9", x"54bb", x"54be", x"54c0", x"54c2", x"54c5", x"54c7", 
    x"54c9", x"54cc", x"54ce", x"54d0", x"54d3", x"54d5", x"54d7", x"54da", 
    x"54dc", x"54df", x"54e1", x"54e3", x"54e6", x"54e8", x"54ea", x"54ed", 
    x"54ef", x"54f1", x"54f4", x"54f6", x"54f8", x"54fb", x"54fd", x"54ff", 
    x"5502", x"5504", x"5506", x"5509", x"550b", x"550e", x"5510", x"5512", 
    x"5515", x"5517", x"5519", x"551c", x"551e", x"5520", x"5523", x"5525", 
    x"5527", x"552a", x"552c", x"552e", x"5531", x"5533", x"5535", x"5538", 
    x"553a", x"553c", x"553f", x"5541", x"5543", x"5546", x"5548", x"554b", 
    x"554d", x"554f", x"5552", x"5554", x"5556", x"5559", x"555b", x"555d", 
    x"5560", x"5562", x"5564", x"5567", x"5569", x"556b", x"556e", x"5570", 
    x"5572", x"5575", x"5577", x"5579", x"557c", x"557e", x"5580", x"5583", 
    x"5585", x"5587", x"558a", x"558c", x"558e", x"5591", x"5593", x"5595", 
    x"5598", x"559a", x"559c", x"559f", x"55a1", x"55a3", x"55a6", x"55a8", 
    x"55aa", x"55ad", x"55af", x"55b1", x"55b4", x"55b6", x"55b8", x"55bb", 
    x"55bd", x"55bf", x"55c2", x"55c4", x"55c6", x"55c9", x"55cb", x"55cd", 
    x"55d0", x"55d2", x"55d4", x"55d7", x"55d9", x"55db", x"55de", x"55e0", 
    x"55e2", x"55e5", x"55e7", x"55e9", x"55ec", x"55ee", x"55f0", x"55f3", 
    x"55f5", x"55f7", x"55fa", x"55fc", x"55fe", x"5601", x"5603", x"5605", 
    x"5608", x"560a", x"560c", x"560f", x"5611", x"5613", x"5616", x"5618", 
    x"561a", x"561d", x"561f", x"5621", x"5623", x"5626", x"5628", x"562a", 
    x"562d", x"562f", x"5631", x"5634", x"5636", x"5638", x"563b", x"563d", 
    x"563f", x"5642", x"5644", x"5646", x"5649", x"564b", x"564d", x"5650", 
    x"5652", x"5654", x"5657", x"5659", x"565b", x"565e", x"5660", x"5662", 
    x"5664", x"5667", x"5669", x"566b", x"566e", x"5670", x"5672", x"5675", 
    x"5677", x"5679", x"567c", x"567e", x"5680", x"5683", x"5685", x"5687", 
    x"568a", x"568c", x"568e", x"5690", x"5693", x"5695", x"5697", x"569a", 
    x"569c", x"569e", x"56a1", x"56a3", x"56a5", x"56a8", x"56aa", x"56ac", 
    x"56af", x"56b1", x"56b3", x"56b5", x"56b8", x"56ba", x"56bc", x"56bf", 
    x"56c1", x"56c3", x"56c6", x"56c8", x"56ca", x"56cd", x"56cf", x"56d1", 
    x"56d3", x"56d6", x"56d8", x"56da", x"56dd", x"56df", x"56e1", x"56e4", 
    x"56e6", x"56e8", x"56eb", x"56ed", x"56ef", x"56f1", x"56f4", x"56f6", 
    x"56f8", x"56fb", x"56fd", x"56ff", x"5702", x"5704", x"5706", x"5709", 
    x"570b", x"570d", x"570f", x"5712", x"5714", x"5716", x"5719", x"571b", 
    x"571d", x"5720", x"5722", x"5724", x"5726", x"5729", x"572b", x"572d", 
    x"5730", x"5732", x"5734", x"5737", x"5739", x"573b", x"573d", x"5740", 
    x"5742", x"5744", x"5747", x"5749", x"574b", x"574e", x"5750", x"5752", 
    x"5754", x"5757", x"5759", x"575b", x"575e", x"5760", x"5762", x"5765", 
    x"5767", x"5769", x"576b", x"576e", x"5770", x"5772", x"5775", x"5777", 
    x"5779", x"577b", x"577e", x"5780", x"5782", x"5785", x"5787", x"5789", 
    x"578b", x"578e", x"5790", x"5792", x"5795", x"5797", x"5799", x"579c", 
    x"579e", x"57a0", x"57a2", x"57a5", x"57a7", x"57a9", x"57ac", x"57ae", 
    x"57b0", x"57b2", x"57b5", x"57b7", x"57b9", x"57bc", x"57be", x"57c0", 
    x"57c2", x"57c5", x"57c7", x"57c9", x"57cc", x"57ce", x"57d0", x"57d2", 
    x"57d5", x"57d7", x"57d9", x"57dc", x"57de", x"57e0", x"57e2", x"57e5", 
    x"57e7", x"57e9", x"57ec", x"57ee", x"57f0", x"57f2", x"57f5", x"57f7", 
    x"57f9", x"57fc", x"57fe", x"5800", x"5802", x"5805", x"5807", x"5809", 
    x"580c", x"580e", x"5810", x"5812", x"5815", x"5817", x"5819", x"581b", 
    x"581e", x"5820", x"5822", x"5825", x"5827", x"5829", x"582b", x"582e", 
    x"5830", x"5832", x"5835", x"5837", x"5839", x"583b", x"583e", x"5840", 
    x"5842", x"5844", x"5847", x"5849", x"584b", x"584e", x"5850", x"5852", 
    x"5854", x"5857", x"5859", x"585b", x"585d", x"5860", x"5862", x"5864", 
    x"5867", x"5869", x"586b", x"586d", x"5870", x"5872", x"5874", x"5876", 
    x"5879", x"587b", x"587d", x"5880", x"5882", x"5884", x"5886", x"5889", 
    x"588b", x"588d", x"588f", x"5892", x"5894", x"5896", x"5898", x"589b", 
    x"589d", x"589f", x"58a2", x"58a4", x"58a6", x"58a8", x"58ab", x"58ad", 
    x"58af", x"58b1", x"58b4", x"58b6", x"58b8", x"58ba", x"58bd", x"58bf", 
    x"58c1", x"58c4", x"58c6", x"58c8", x"58ca", x"58cd", x"58cf", x"58d1", 
    x"58d3", x"58d6", x"58d8", x"58da", x"58dc", x"58df", x"58e1", x"58e3", 
    x"58e5", x"58e8", x"58ea", x"58ec", x"58ee", x"58f1", x"58f3", x"58f5", 
    x"58f8", x"58fa", x"58fc", x"58fe", x"5901", x"5903", x"5905", x"5907", 
    x"590a", x"590c", x"590e", x"5910", x"5913", x"5915", x"5917", x"5919", 
    x"591c", x"591e", x"5920", x"5922", x"5925", x"5927", x"5929", x"592b", 
    x"592e", x"5930", x"5932", x"5934", x"5937", x"5939", x"593b", x"593d", 
    x"5940", x"5942", x"5944", x"5946", x"5949", x"594b", x"594d", x"594f", 
    x"5952", x"5954", x"5956", x"5958", x"595b", x"595d", x"595f", x"5961", 
    x"5964", x"5966", x"5968", x"596a", x"596d", x"596f", x"5971", x"5973", 
    x"5976", x"5978", x"597a", x"597c", x"597f", x"5981", x"5983", x"5985", 
    x"5988", x"598a", x"598c", x"598e", x"5991", x"5993", x"5995", x"5997", 
    x"599a", x"599c", x"599e", x"59a0", x"59a3", x"59a5", x"59a7", x"59a9", 
    x"59ac", x"59ae", x"59b0", x"59b2", x"59b5", x"59b7", x"59b9", x"59bb", 
    x"59bd", x"59c0", x"59c2", x"59c4", x"59c6", x"59c9", x"59cb", x"59cd", 
    x"59cf", x"59d2", x"59d4", x"59d6", x"59d8", x"59db", x"59dd", x"59df", 
    x"59e1", x"59e4", x"59e6", x"59e8", x"59ea", x"59ec", x"59ef", x"59f1", 
    x"59f3", x"59f5", x"59f8", x"59fa", x"59fc", x"59fe", x"5a01", x"5a03", 
    x"5a05", x"5a07", x"5a0a", x"5a0c", x"5a0e", x"5a10", x"5a12", x"5a15", 
    x"5a17", x"5a19", x"5a1b", x"5a1e", x"5a20", x"5a22", x"5a24", x"5a27", 
    x"5a29", x"5a2b", x"5a2d", x"5a2f", x"5a32", x"5a34", x"5a36", x"5a38", 
    x"5a3b", x"5a3d", x"5a3f", x"5a41", x"5a43", x"5a46", x"5a48", x"5a4a", 
    x"5a4c", x"5a4f", x"5a51", x"5a53", x"5a55", x"5a58", x"5a5a", x"5a5c", 
    x"5a5e", x"5a60", x"5a63", x"5a65", x"5a67", x"5a69", x"5a6c", x"5a6e", 
    x"5a70", x"5a72", x"5a74", x"5a77", x"5a79", x"5a7b", x"5a7d", x"5a80", 
    x"5a82", x"5a84", x"5a86", x"5a88", x"5a8b", x"5a8d", x"5a8f", x"5a91", 
    x"5a94", x"5a96", x"5a98", x"5a9a", x"5a9c", x"5a9f", x"5aa1", x"5aa3", 
    x"5aa5", x"5aa8", x"5aaa", x"5aac", x"5aae", x"5ab0", x"5ab3", x"5ab5", 
    x"5ab7", x"5ab9", x"5abb", x"5abe", x"5ac0", x"5ac2", x"5ac4", x"5ac7", 
    x"5ac9", x"5acb", x"5acd", x"5acf", x"5ad2", x"5ad4", x"5ad6", x"5ad8", 
    x"5ada", x"5add", x"5adf", x"5ae1", x"5ae3", x"5ae6", x"5ae8", x"5aea", 
    x"5aec", x"5aee", x"5af1", x"5af3", x"5af5", x"5af7", x"5af9", x"5afc", 
    x"5afe", x"5b00", x"5b02", x"5b04", x"5b07", x"5b09", x"5b0b", x"5b0d", 
    x"5b0f", x"5b12", x"5b14", x"5b16", x"5b18", x"5b1b", x"5b1d", x"5b1f", 
    x"5b21", x"5b23", x"5b26", x"5b28", x"5b2a", x"5b2c", x"5b2e", x"5b31", 
    x"5b33", x"5b35", x"5b37", x"5b39", x"5b3c", x"5b3e", x"5b40", x"5b42", 
    x"5b44", x"5b47", x"5b49", x"5b4b", x"5b4d", x"5b4f", x"5b52", x"5b54", 
    x"5b56", x"5b58", x"5b5a", x"5b5d", x"5b5f", x"5b61", x"5b63", x"5b65", 
    x"5b68", x"5b6a", x"5b6c", x"5b6e", x"5b70", x"5b73", x"5b75", x"5b77", 
    x"5b79", x"5b7b", x"5b7e", x"5b80", x"5b82", x"5b84", x"5b86", x"5b89", 
    x"5b8b", x"5b8d", x"5b8f", x"5b91", x"5b94", x"5b96", x"5b98", x"5b9a", 
    x"5b9c", x"5b9f", x"5ba1", x"5ba3", x"5ba5", x"5ba7", x"5baa", x"5bac", 
    x"5bae", x"5bb0", x"5bb2", x"5bb4", x"5bb7", x"5bb9", x"5bbb", x"5bbd", 
    x"5bbf", x"5bc2", x"5bc4", x"5bc6", x"5bc8", x"5bca", x"5bcd", x"5bcf", 
    x"5bd1", x"5bd3", x"5bd5", x"5bd8", x"5bda", x"5bdc", x"5bde", x"5be0", 
    x"5be2", x"5be5", x"5be7", x"5be9", x"5beb", x"5bed", x"5bf0", x"5bf2", 
    x"5bf4", x"5bf6", x"5bf8", x"5bfa", x"5bfd", x"5bff", x"5c01", x"5c03", 
    x"5c05", x"5c08", x"5c0a", x"5c0c", x"5c0e", x"5c10", x"5c13", x"5c15", 
    x"5c17", x"5c19", x"5c1b", x"5c1d", x"5c20", x"5c22", x"5c24", x"5c26", 
    x"5c28", x"5c2b", x"5c2d", x"5c2f", x"5c31", x"5c33", x"5c35", x"5c38", 
    x"5c3a", x"5c3c", x"5c3e", x"5c40", x"5c42", x"5c45", x"5c47", x"5c49", 
    x"5c4b", x"5c4d", x"5c50", x"5c52", x"5c54", x"5c56", x"5c58", x"5c5a", 
    x"5c5d", x"5c5f", x"5c61", x"5c63", x"5c65", x"5c67", x"5c6a", x"5c6c", 
    x"5c6e", x"5c70", x"5c72", x"5c74", x"5c77", x"5c79", x"5c7b", x"5c7d", 
    x"5c7f", x"5c82", x"5c84", x"5c86", x"5c88", x"5c8a", x"5c8c", x"5c8f", 
    x"5c91", x"5c93", x"5c95", x"5c97", x"5c99", x"5c9c", x"5c9e", x"5ca0", 
    x"5ca2", x"5ca4", x"5ca6", x"5ca9", x"5cab", x"5cad", x"5caf", x"5cb1", 
    x"5cb3", x"5cb6", x"5cb8", x"5cba", x"5cbc", x"5cbe", x"5cc0", x"5cc3", 
    x"5cc5", x"5cc7", x"5cc9", x"5ccb", x"5ccd", x"5cd0", x"5cd2", x"5cd4", 
    x"5cd6", x"5cd8", x"5cda", x"5cdd", x"5cdf", x"5ce1", x"5ce3", x"5ce5", 
    x"5ce7", x"5ce9", x"5cec", x"5cee", x"5cf0", x"5cf2", x"5cf4", x"5cf6", 
    x"5cf9", x"5cfb", x"5cfd", x"5cff", x"5d01", x"5d03", x"5d06", x"5d08", 
    x"5d0a", x"5d0c", x"5d0e", x"5d10", x"5d13", x"5d15", x"5d17", x"5d19", 
    x"5d1b", x"5d1d", x"5d1f", x"5d22", x"5d24", x"5d26", x"5d28", x"5d2a", 
    x"5d2c", x"5d2f", x"5d31", x"5d33", x"5d35", x"5d37", x"5d39", x"5d3b", 
    x"5d3e", x"5d40", x"5d42", x"5d44", x"5d46", x"5d48", x"5d4b", x"5d4d", 
    x"5d4f", x"5d51", x"5d53", x"5d55", x"5d57", x"5d5a", x"5d5c", x"5d5e", 
    x"5d60", x"5d62", x"5d64", x"5d66", x"5d69", x"5d6b", x"5d6d", x"5d6f", 
    x"5d71", x"5d73", x"5d75", x"5d78", x"5d7a", x"5d7c", x"5d7e", x"5d80", 
    x"5d82", x"5d84", x"5d87", x"5d89", x"5d8b", x"5d8d", x"5d8f", x"5d91", 
    x"5d94", x"5d96", x"5d98", x"5d9a", x"5d9c", x"5d9e", x"5da0", x"5da3", 
    x"5da5", x"5da7", x"5da9", x"5dab", x"5dad", x"5daf", x"5db1", x"5db4", 
    x"5db6", x"5db8", x"5dba", x"5dbc", x"5dbe", x"5dc0", x"5dc3", x"5dc5", 
    x"5dc7", x"5dc9", x"5dcb", x"5dcd", x"5dcf", x"5dd2", x"5dd4", x"5dd6", 
    x"5dd8", x"5dda", x"5ddc", x"5dde", x"5de1", x"5de3", x"5de5", x"5de7", 
    x"5de9", x"5deb", x"5ded", x"5def", x"5df2", x"5df4", x"5df6", x"5df8", 
    x"5dfa", x"5dfc", x"5dfe", x"5e01", x"5e03", x"5e05", x"5e07", x"5e09", 
    x"5e0b", x"5e0d", x"5e0f", x"5e12", x"5e14", x"5e16", x"5e18", x"5e1a", 
    x"5e1c", x"5e1e", x"5e20", x"5e23", x"5e25", x"5e27", x"5e29", x"5e2b", 
    x"5e2d", x"5e2f", x"5e32", x"5e34", x"5e36", x"5e38", x"5e3a", x"5e3c", 
    x"5e3e", x"5e40", x"5e43", x"5e45", x"5e47", x"5e49", x"5e4b", x"5e4d", 
    x"5e4f", x"5e51", x"5e54", x"5e56", x"5e58", x"5e5a", x"5e5c", x"5e5e", 
    x"5e60", x"5e62", x"5e64", x"5e67", x"5e69", x"5e6b", x"5e6d", x"5e6f", 
    x"5e71", x"5e73", x"5e75", x"5e78", x"5e7a", x"5e7c", x"5e7e", x"5e80", 
    x"5e82", x"5e84", x"5e86", x"5e89", x"5e8b", x"5e8d", x"5e8f", x"5e91", 
    x"5e93", x"5e95", x"5e97", x"5e99", x"5e9c", x"5e9e", x"5ea0", x"5ea2", 
    x"5ea4", x"5ea6", x"5ea8", x"5eaa", x"5ead", x"5eaf", x"5eb1", x"5eb3", 
    x"5eb5", x"5eb7", x"5eb9", x"5ebb", x"5ebd", x"5ec0", x"5ec2", x"5ec4", 
    x"5ec6", x"5ec8", x"5eca", x"5ecc", x"5ece", x"5ed0", x"5ed3", x"5ed5", 
    x"5ed7", x"5ed9", x"5edb", x"5edd", x"5edf", x"5ee1", x"5ee3", x"5ee6", 
    x"5ee8", x"5eea", x"5eec", x"5eee", x"5ef0", x"5ef2", x"5ef4", x"5ef6", 
    x"5ef8", x"5efb", x"5efd", x"5eff", x"5f01", x"5f03", x"5f05", x"5f07", 
    x"5f09", x"5f0b", x"5f0e", x"5f10", x"5f12", x"5f14", x"5f16", x"5f18", 
    x"5f1a", x"5f1c", x"5f1e", x"5f20", x"5f23", x"5f25", x"5f27", x"5f29", 
    x"5f2b", x"5f2d", x"5f2f", x"5f31", x"5f33", x"5f35", x"5f38", x"5f3a", 
    x"5f3c", x"5f3e", x"5f40", x"5f42", x"5f44", x"5f46", x"5f48", x"5f4a", 
    x"5f4d", x"5f4f", x"5f51", x"5f53", x"5f55", x"5f57", x"5f59", x"5f5b", 
    x"5f5d", x"5f5f", x"5f61", x"5f64", x"5f66", x"5f68", x"5f6a", x"5f6c", 
    x"5f6e", x"5f70", x"5f72", x"5f74", x"5f76", x"5f79", x"5f7b", x"5f7d", 
    x"5f7f", x"5f81", x"5f83", x"5f85", x"5f87", x"5f89", x"5f8b", x"5f8d", 
    x"5f90", x"5f92", x"5f94", x"5f96", x"5f98", x"5f9a", x"5f9c", x"5f9e", 
    x"5fa0", x"5fa2", x"5fa4", x"5fa7", x"5fa9", x"5fab", x"5fad", x"5faf", 
    x"5fb1", x"5fb3", x"5fb5", x"5fb7", x"5fb9", x"5fbb", x"5fbd", x"5fc0", 
    x"5fc2", x"5fc4", x"5fc6", x"5fc8", x"5fca", x"5fcc", x"5fce", x"5fd0", 
    x"5fd2", x"5fd4", x"5fd6", x"5fd9", x"5fdb", x"5fdd", x"5fdf", x"5fe1", 
    x"5fe3", x"5fe5", x"5fe7", x"5fe9", x"5feb", x"5fed", x"5fef", x"5ff2", 
    x"5ff4", x"5ff6", x"5ff8", x"5ffa", x"5ffc", x"5ffe", x"6000", x"6002", 
    x"6004", x"6006", x"6008", x"600a", x"600d", x"600f", x"6011", x"6013", 
    x"6015", x"6017", x"6019", x"601b", x"601d", x"601f", x"6021", x"6023", 
    x"6025", x"6028", x"602a", x"602c", x"602e", x"6030", x"6032", x"6034", 
    x"6036", x"6038", x"603a", x"603c", x"603e", x"6040", x"6042", x"6045", 
    x"6047", x"6049", x"604b", x"604d", x"604f", x"6051", x"6053", x"6055", 
    x"6057", x"6059", x"605b", x"605d", x"605f", x"6061", x"6064", x"6066", 
    x"6068", x"606a", x"606c", x"606e", x"6070", x"6072", x"6074", x"6076", 
    x"6078", x"607a", x"607c", x"607e", x"6080", x"6083", x"6085", x"6087", 
    x"6089", x"608b", x"608d", x"608f", x"6091", x"6093", x"6095", x"6097", 
    x"6099", x"609b", x"609d", x"609f", x"60a1", x"60a4", x"60a6", x"60a8", 
    x"60aa", x"60ac", x"60ae", x"60b0", x"60b2", x"60b4", x"60b6", x"60b8", 
    x"60ba", x"60bc", x"60be", x"60c0", x"60c2", x"60c4", x"60c6", x"60c9", 
    x"60cb", x"60cd", x"60cf", x"60d1", x"60d3", x"60d5", x"60d7", x"60d9", 
    x"60db", x"60dd", x"60df", x"60e1", x"60e3", x"60e5", x"60e7", x"60e9", 
    x"60eb", x"60ee", x"60f0", x"60f2", x"60f4", x"60f6", x"60f8", x"60fa", 
    x"60fc", x"60fe", x"6100", x"6102", x"6104", x"6106", x"6108", x"610a", 
    x"610c", x"610e", x"6110", x"6112", x"6114", x"6117", x"6119", x"611b", 
    x"611d", x"611f", x"6121", x"6123", x"6125", x"6127", x"6129", x"612b", 
    x"612d", x"612f", x"6131", x"6133", x"6135", x"6137", x"6139", x"613b", 
    x"613d", x"613f", x"6141", x"6143", x"6146", x"6148", x"614a", x"614c", 
    x"614e", x"6150", x"6152", x"6154", x"6156", x"6158", x"615a", x"615c", 
    x"615e", x"6160", x"6162", x"6164", x"6166", x"6168", x"616a", x"616c", 
    x"616e", x"6170", x"6172", x"6174", x"6176", x"6179", x"617b", x"617d", 
    x"617f", x"6181", x"6183", x"6185", x"6187", x"6189", x"618b", x"618d", 
    x"618f", x"6191", x"6193", x"6195", x"6197", x"6199", x"619b", x"619d", 
    x"619f", x"61a1", x"61a3", x"61a5", x"61a7", x"61a9", x"61ab", x"61ad", 
    x"61af", x"61b1", x"61b3", x"61b5", x"61b8", x"61ba", x"61bc", x"61be", 
    x"61c0", x"61c2", x"61c4", x"61c6", x"61c8", x"61ca", x"61cc", x"61ce", 
    x"61d0", x"61d2", x"61d4", x"61d6", x"61d8", x"61da", x"61dc", x"61de", 
    x"61e0", x"61e2", x"61e4", x"61e6", x"61e8", x"61ea", x"61ec", x"61ee", 
    x"61f0", x"61f2", x"61f4", x"61f6", x"61f8", x"61fa", x"61fc", x"61fe", 
    x"6200", x"6202", x"6204", x"6206", x"6208", x"620b", x"620d", x"620f", 
    x"6211", x"6213", x"6215", x"6217", x"6219", x"621b", x"621d", x"621f", 
    x"6221", x"6223", x"6225", x"6227", x"6229", x"622b", x"622d", x"622f", 
    x"6231", x"6233", x"6235", x"6237", x"6239", x"623b", x"623d", x"623f", 
    x"6241", x"6243", x"6245", x"6247", x"6249", x"624b", x"624d", x"624f", 
    x"6251", x"6253", x"6255", x"6257", x"6259", x"625b", x"625d", x"625f", 
    x"6261", x"6263", x"6265", x"6267", x"6269", x"626b", x"626d", x"626f", 
    x"6271", x"6273", x"6275", x"6277", x"6279", x"627b", x"627d", x"627f", 
    x"6281", x"6283", x"6285", x"6287", x"6289", x"628b", x"628d", x"628f", 
    x"6291", x"6293", x"6295", x"6297", x"6299", x"629b", x"629d", x"629f", 
    x"62a1", x"62a3", x"62a5", x"62a7", x"62a9", x"62ab", x"62ad", x"62af", 
    x"62b1", x"62b3", x"62b5", x"62b7", x"62b9", x"62bb", x"62bd", x"62bf", 
    x"62c1", x"62c3", x"62c5", x"62c7", x"62c9", x"62cb", x"62cd", x"62cf", 
    x"62d1", x"62d3", x"62d5", x"62d7", x"62d9", x"62db", x"62dd", x"62df", 
    x"62e1", x"62e3", x"62e5", x"62e7", x"62e9", x"62eb", x"62ed", x"62ef", 
    x"62f1", x"62f3", x"62f5", x"62f7", x"62f9", x"62fb", x"62fd", x"62ff", 
    x"6301", x"6303", x"6305", x"6307", x"6309", x"630b", x"630d", x"630f", 
    x"6311", x"6313", x"6315", x"6317", x"6319", x"631b", x"631d", x"631f", 
    x"6321", x"6323", x"6325", x"6327", x"6329", x"632b", x"632d", x"632f", 
    x"6331", x"6333", x"6335", x"6337", x"6339", x"633b", x"633d", x"633f", 
    x"6341", x"6343", x"6345", x"6347", x"6349", x"634b", x"634d", x"634f", 
    x"6351", x"6353", x"6355", x"6357", x"6359", x"635b", x"635d", x"635e", 
    x"6360", x"6362", x"6364", x"6366", x"6368", x"636a", x"636c", x"636e", 
    x"6370", x"6372", x"6374", x"6376", x"6378", x"637a", x"637c", x"637e", 
    x"6380", x"6382", x"6384", x"6386", x"6388", x"638a", x"638c", x"638e", 
    x"6390", x"6392", x"6394", x"6396", x"6398", x"639a", x"639c", x"639e", 
    x"63a0", x"63a2", x"63a4", x"63a6", x"63a8", x"63aa", x"63ac", x"63ae", 
    x"63af", x"63b1", x"63b3", x"63b5", x"63b7", x"63b9", x"63bb", x"63bd", 
    x"63bf", x"63c1", x"63c3", x"63c5", x"63c7", x"63c9", x"63cb", x"63cd", 
    x"63cf", x"63d1", x"63d3", x"63d5", x"63d7", x"63d9", x"63db", x"63dd", 
    x"63df", x"63e1", x"63e3", x"63e5", x"63e7", x"63e9", x"63ea", x"63ec", 
    x"63ee", x"63f0", x"63f2", x"63f4", x"63f6", x"63f8", x"63fa", x"63fc", 
    x"63fe", x"6400", x"6402", x"6404", x"6406", x"6408", x"640a", x"640c", 
    x"640e", x"6410", x"6412", x"6414", x"6416", x"6418", x"641a", x"641c", 
    x"641d", x"641f", x"6421", x"6423", x"6425", x"6427", x"6429", x"642b", 
    x"642d", x"642f", x"6431", x"6433", x"6435", x"6437", x"6439", x"643b", 
    x"643d", x"643f", x"6441", x"6443", x"6445", x"6447", x"6448", x"644a", 
    x"644c", x"644e", x"6450", x"6452", x"6454", x"6456", x"6458", x"645a", 
    x"645c", x"645e", x"6460", x"6462", x"6464", x"6466", x"6468", x"646a", 
    x"646c", x"646e", x"646f", x"6471", x"6473", x"6475", x"6477", x"6479", 
    x"647b", x"647d", x"647f", x"6481", x"6483", x"6485", x"6487", x"6489", 
    x"648b", x"648d", x"648f", x"6491", x"6492", x"6494", x"6496", x"6498", 
    x"649a", x"649c", x"649e", x"64a0", x"64a2", x"64a4", x"64a6", x"64a8", 
    x"64aa", x"64ac", x"64ae", x"64b0", x"64b2", x"64b3", x"64b5", x"64b7", 
    x"64b9", x"64bb", x"64bd", x"64bf", x"64c1", x"64c3", x"64c5", x"64c7", 
    x"64c9", x"64cb", x"64cd", x"64cf", x"64d1", x"64d2", x"64d4", x"64d6", 
    x"64d8", x"64da", x"64dc", x"64de", x"64e0", x"64e2", x"64e4", x"64e6", 
    x"64e8", x"64ea", x"64ec", x"64ee", x"64ef", x"64f1", x"64f3", x"64f5", 
    x"64f7", x"64f9", x"64fb", x"64fd", x"64ff", x"6501", x"6503", x"6505", 
    x"6507", x"6509", x"650a", x"650c", x"650e", x"6510", x"6512", x"6514", 
    x"6516", x"6518", x"651a", x"651c", x"651e", x"6520", x"6522", x"6524", 
    x"6525", x"6527", x"6529", x"652b", x"652d", x"652f", x"6531", x"6533", 
    x"6535", x"6537", x"6539", x"653b", x"653d", x"653e", x"6540", x"6542", 
    x"6544", x"6546", x"6548", x"654a", x"654c", x"654e", x"6550", x"6552", 
    x"6554", x"6556", x"6557", x"6559", x"655b", x"655d", x"655f", x"6561", 
    x"6563", x"6565", x"6567", x"6569", x"656b", x"656d", x"656e", x"6570", 
    x"6572", x"6574", x"6576", x"6578", x"657a", x"657c", x"657e", x"6580", 
    x"6582", x"6584", x"6585", x"6587", x"6589", x"658b", x"658d", x"658f", 
    x"6591", x"6593", x"6595", x"6597", x"6599", x"659a", x"659c", x"659e", 
    x"65a0", x"65a2", x"65a4", x"65a6", x"65a8", x"65aa", x"65ac", x"65ae", 
    x"65af", x"65b1", x"65b3", x"65b5", x"65b7", x"65b9", x"65bb", x"65bd", 
    x"65bf", x"65c1", x"65c3", x"65c4", x"65c6", x"65c8", x"65ca", x"65cc", 
    x"65ce", x"65d0", x"65d2", x"65d4", x"65d6", x"65d7", x"65d9", x"65db", 
    x"65dd", x"65df", x"65e1", x"65e3", x"65e5", x"65e7", x"65e9", x"65ea", 
    x"65ec", x"65ee", x"65f0", x"65f2", x"65f4", x"65f6", x"65f8", x"65fa", 
    x"65fc", x"65fd", x"65ff", x"6601", x"6603", x"6605", x"6607", x"6609", 
    x"660b", x"660d", x"660f", x"6610", x"6612", x"6614", x"6616", x"6618", 
    x"661a", x"661c", x"661e", x"6620", x"6622", x"6623", x"6625", x"6627", 
    x"6629", x"662b", x"662d", x"662f", x"6631", x"6633", x"6634", x"6636", 
    x"6638", x"663a", x"663c", x"663e", x"6640", x"6642", x"6644", x"6645", 
    x"6647", x"6649", x"664b", x"664d", x"664f", x"6651", x"6653", x"6655", 
    x"6656", x"6658", x"665a", x"665c", x"665e", x"6660", x"6662", x"6664", 
    x"6666", x"6667", x"6669", x"666b", x"666d", x"666f", x"6671", x"6673", 
    x"6675", x"6676", x"6678", x"667a", x"667c", x"667e", x"6680", x"6682", 
    x"6684", x"6686", x"6687", x"6689", x"668b", x"668d", x"668f", x"6691", 
    x"6693", x"6695", x"6696", x"6698", x"669a", x"669c", x"669e", x"66a0", 
    x"66a2", x"66a4", x"66a5", x"66a7", x"66a9", x"66ab", x"66ad", x"66af", 
    x"66b1", x"66b3", x"66b4", x"66b6", x"66b8", x"66ba", x"66bc", x"66be", 
    x"66c0", x"66c2", x"66c3", x"66c5", x"66c7", x"66c9", x"66cb", x"66cd", 
    x"66cf", x"66d1", x"66d2", x"66d4", x"66d6", x"66d8", x"66da", x"66dc", 
    x"66de", x"66e0", x"66e1", x"66e3", x"66e5", x"66e7", x"66e9", x"66eb", 
    x"66ed", x"66ee", x"66f0", x"66f2", x"66f4", x"66f6", x"66f8", x"66fa", 
    x"66fc", x"66fd", x"66ff", x"6701", x"6703", x"6705", x"6707", x"6709", 
    x"670a", x"670c", x"670e", x"6710", x"6712", x"6714", x"6716", x"6718", 
    x"6719", x"671b", x"671d", x"671f", x"6721", x"6723", x"6725", x"6726", 
    x"6728", x"672a", x"672c", x"672e", x"6730", x"6732", x"6733", x"6735", 
    x"6737", x"6739", x"673b", x"673d", x"673f", x"6740", x"6742", x"6744", 
    x"6746", x"6748", x"674a", x"674c", x"674d", x"674f", x"6751", x"6753", 
    x"6755", x"6757", x"6759", x"675a", x"675c", x"675e", x"6760", x"6762", 
    x"6764", x"6765", x"6767", x"6769", x"676b", x"676d", x"676f", x"6771", 
    x"6772", x"6774", x"6776", x"6778", x"677a", x"677c", x"677e", x"677f", 
    x"6781", x"6783", x"6785", x"6787", x"6789", x"678a", x"678c", x"678e", 
    x"6790", x"6792", x"6794", x"6796", x"6797", x"6799", x"679b", x"679d", 
    x"679f", x"67a1", x"67a2", x"67a4", x"67a6", x"67a8", x"67aa", x"67ac", 
    x"67ae", x"67af", x"67b1", x"67b3", x"67b5", x"67b7", x"67b9", x"67ba", 
    x"67bc", x"67be", x"67c0", x"67c2", x"67c4", x"67c5", x"67c7", x"67c9", 
    x"67cb", x"67cd", x"67cf", x"67d0", x"67d2", x"67d4", x"67d6", x"67d8", 
    x"67da", x"67dc", x"67dd", x"67df", x"67e1", x"67e3", x"67e5", x"67e7", 
    x"67e8", x"67ea", x"67ec", x"67ee", x"67f0", x"67f2", x"67f3", x"67f5", 
    x"67f7", x"67f9", x"67fb", x"67fd", x"67fe", x"6800", x"6802", x"6804", 
    x"6806", x"6807", x"6809", x"680b", x"680d", x"680f", x"6811", x"6812", 
    x"6814", x"6816", x"6818", x"681a", x"681c", x"681d", x"681f", x"6821", 
    x"6823", x"6825", x"6827", x"6828", x"682a", x"682c", x"682e", x"6830", 
    x"6832", x"6833", x"6835", x"6837", x"6839", x"683b", x"683c", x"683e", 
    x"6840", x"6842", x"6844", x"6846", x"6847", x"6849", x"684b", x"684d", 
    x"684f", x"6851", x"6852", x"6854", x"6856", x"6858", x"685a", x"685b", 
    x"685d", x"685f", x"6861", x"6863", x"6865", x"6866", x"6868", x"686a", 
    x"686c", x"686e", x"686f", x"6871", x"6873", x"6875", x"6877", x"6879", 
    x"687a", x"687c", x"687e", x"6880", x"6882", x"6883", x"6885", x"6887", 
    x"6889", x"688b", x"688c", x"688e", x"6890", x"6892", x"6894", x"6896", 
    x"6897", x"6899", x"689b", x"689d", x"689f", x"68a0", x"68a2", x"68a4", 
    x"68a6", x"68a8", x"68a9", x"68ab", x"68ad", x"68af", x"68b1", x"68b2", 
    x"68b4", x"68b6", x"68b8", x"68ba", x"68bb", x"68bd", x"68bf", x"68c1", 
    x"68c3", x"68c5", x"68c6", x"68c8", x"68ca", x"68cc", x"68ce", x"68cf", 
    x"68d1", x"68d3", x"68d5", x"68d7", x"68d8", x"68da", x"68dc", x"68de", 
    x"68e0", x"68e1", x"68e3", x"68e5", x"68e7", x"68e9", x"68ea", x"68ec", 
    x"68ee", x"68f0", x"68f2", x"68f3", x"68f5", x"68f7", x"68f9", x"68fb", 
    x"68fc", x"68fe", x"6900", x"6902", x"6904", x"6905", x"6907", x"6909", 
    x"690b", x"690d", x"690e", x"6910", x"6912", x"6914", x"6915", x"6917", 
    x"6919", x"691b", x"691d", x"691e", x"6920", x"6922", x"6924", x"6926", 
    x"6927", x"6929", x"692b", x"692d", x"692f", x"6930", x"6932", x"6934", 
    x"6936", x"6938", x"6939", x"693b", x"693d", x"693f", x"6940", x"6942", 
    x"6944", x"6946", x"6948", x"6949", x"694b", x"694d", x"694f", x"6951", 
    x"6952", x"6954", x"6956", x"6958", x"6959", x"695b", x"695d", x"695f", 
    x"6961", x"6962", x"6964", x"6966", x"6968", x"696a", x"696b", x"696d", 
    x"696f", x"6971", x"6972", x"6974", x"6976", x"6978", x"697a", x"697b", 
    x"697d", x"697f", x"6981", x"6982", x"6984", x"6986", x"6988", x"698a", 
    x"698b", x"698d", x"698f", x"6991", x"6992", x"6994", x"6996", x"6998", 
    x"699a", x"699b", x"699d", x"699f", x"69a1", x"69a2", x"69a4", x"69a6", 
    x"69a8", x"69a9", x"69ab", x"69ad", x"69af", x"69b1", x"69b2", x"69b4", 
    x"69b6", x"69b8", x"69b9", x"69bb", x"69bd", x"69bf", x"69c1", x"69c2", 
    x"69c4", x"69c6", x"69c8", x"69c9", x"69cb", x"69cd", x"69cf", x"69d0", 
    x"69d2", x"69d4", x"69d6", x"69d8", x"69d9", x"69db", x"69dd", x"69df", 
    x"69e0", x"69e2", x"69e4", x"69e6", x"69e7", x"69e9", x"69eb", x"69ed", 
    x"69ee", x"69f0", x"69f2", x"69f4", x"69f6", x"69f7", x"69f9", x"69fb", 
    x"69fd", x"69fe", x"6a00", x"6a02", x"6a04", x"6a05", x"6a07", x"6a09", 
    x"6a0b", x"6a0c", x"6a0e", x"6a10", x"6a12", x"6a13", x"6a15", x"6a17", 
    x"6a19", x"6a1a", x"6a1c", x"6a1e", x"6a20", x"6a21", x"6a23", x"6a25", 
    x"6a27", x"6a29", x"6a2a", x"6a2c", x"6a2e", x"6a30", x"6a31", x"6a33", 
    x"6a35", x"6a37", x"6a38", x"6a3a", x"6a3c", x"6a3e", x"6a3f", x"6a41", 
    x"6a43", x"6a45", x"6a46", x"6a48", x"6a4a", x"6a4c", x"6a4d", x"6a4f", 
    x"6a51", x"6a53", x"6a54", x"6a56", x"6a58", x"6a5a", x"6a5b", x"6a5d", 
    x"6a5f", x"6a61", x"6a62", x"6a64", x"6a66", x"6a68", x"6a69", x"6a6b", 
    x"6a6d", x"6a6f", x"6a70", x"6a72", x"6a74", x"6a75", x"6a77", x"6a79", 
    x"6a7b", x"6a7c", x"6a7e", x"6a80", x"6a82", x"6a83", x"6a85", x"6a87", 
    x"6a89", x"6a8a", x"6a8c", x"6a8e", x"6a90", x"6a91", x"6a93", x"6a95", 
    x"6a97", x"6a98", x"6a9a", x"6a9c", x"6a9e", x"6a9f", x"6aa1", x"6aa3", 
    x"6aa4", x"6aa6", x"6aa8", x"6aaa", x"6aab", x"6aad", x"6aaf", x"6ab1", 
    x"6ab2", x"6ab4", x"6ab6", x"6ab8", x"6ab9", x"6abb", x"6abd", x"6abf", 
    x"6ac0", x"6ac2", x"6ac4", x"6ac5", x"6ac7", x"6ac9", x"6acb", x"6acc", 
    x"6ace", x"6ad0", x"6ad2", x"6ad3", x"6ad5", x"6ad7", x"6ad8", x"6ada", 
    x"6adc", x"6ade", x"6adf", x"6ae1", x"6ae3", x"6ae5", x"6ae6", x"6ae8", 
    x"6aea", x"6aec", x"6aed", x"6aef", x"6af1", x"6af2", x"6af4", x"6af6", 
    x"6af8", x"6af9", x"6afb", x"6afd", x"6afe", x"6b00", x"6b02", x"6b04", 
    x"6b05", x"6b07", x"6b09", x"6b0b", x"6b0c", x"6b0e", x"6b10", x"6b11", 
    x"6b13", x"6b15", x"6b17", x"6b18", x"6b1a", x"6b1c", x"6b1d", x"6b1f", 
    x"6b21", x"6b23", x"6b24", x"6b26", x"6b28", x"6b2a", x"6b2b", x"6b2d", 
    x"6b2f", x"6b30", x"6b32", x"6b34", x"6b36", x"6b37", x"6b39", x"6b3b", 
    x"6b3c", x"6b3e", x"6b40", x"6b42", x"6b43", x"6b45", x"6b47", x"6b48", 
    x"6b4a", x"6b4c", x"6b4e", x"6b4f", x"6b51", x"6b53", x"6b54", x"6b56", 
    x"6b58", x"6b5a", x"6b5b", x"6b5d", x"6b5f", x"6b60", x"6b62", x"6b64", 
    x"6b65", x"6b67", x"6b69", x"6b6b", x"6b6c", x"6b6e", x"6b70", x"6b71", 
    x"6b73", x"6b75", x"6b77", x"6b78", x"6b7a", x"6b7c", x"6b7d", x"6b7f", 
    x"6b81", x"6b83", x"6b84", x"6b86", x"6b88", x"6b89", x"6b8b", x"6b8d", 
    x"6b8e", x"6b90", x"6b92", x"6b94", x"6b95", x"6b97", x"6b99", x"6b9a", 
    x"6b9c", x"6b9e", x"6b9f", x"6ba1", x"6ba3", x"6ba5", x"6ba6", x"6ba8", 
    x"6baa", x"6bab", x"6bad", x"6baf", x"6bb0", x"6bb2", x"6bb4", x"6bb6", 
    x"6bb7", x"6bb9", x"6bbb", x"6bbc", x"6bbe", x"6bc0", x"6bc1", x"6bc3", 
    x"6bc5", x"6bc6", x"6bc8", x"6bca", x"6bcc", x"6bcd", x"6bcf", x"6bd1", 
    x"6bd2", x"6bd4", x"6bd6", x"6bd7", x"6bd9", x"6bdb", x"6bdd", x"6bde", 
    x"6be0", x"6be2", x"6be3", x"6be5", x"6be7", x"6be8", x"6bea", x"6bec", 
    x"6bed", x"6bef", x"6bf1", x"6bf2", x"6bf4", x"6bf6", x"6bf8", x"6bf9", 
    x"6bfb", x"6bfd", x"6bfe", x"6c00", x"6c02", x"6c03", x"6c05", x"6c07", 
    x"6c08", x"6c0a", x"6c0c", x"6c0d", x"6c0f", x"6c11", x"6c12", x"6c14", 
    x"6c16", x"6c18", x"6c19", x"6c1b", x"6c1d", x"6c1e", x"6c20", x"6c22", 
    x"6c23", x"6c25", x"6c27", x"6c28", x"6c2a", x"6c2c", x"6c2d", x"6c2f", 
    x"6c31", x"6c32", x"6c34", x"6c36", x"6c37", x"6c39", x"6c3b", x"6c3c", 
    x"6c3e", x"6c40", x"6c42", x"6c43", x"6c45", x"6c47", x"6c48", x"6c4a", 
    x"6c4c", x"6c4d", x"6c4f", x"6c51", x"6c52", x"6c54", x"6c56", x"6c57", 
    x"6c59", x"6c5b", x"6c5c", x"6c5e", x"6c60", x"6c61", x"6c63", x"6c65", 
    x"6c66", x"6c68", x"6c6a", x"6c6b", x"6c6d", x"6c6f", x"6c70", x"6c72", 
    x"6c74", x"6c75", x"6c77", x"6c79", x"6c7a", x"6c7c", x"6c7e", x"6c7f", 
    x"6c81", x"6c83", x"6c84", x"6c86", x"6c88", x"6c89", x"6c8b", x"6c8d", 
    x"6c8e", x"6c90", x"6c92", x"6c93", x"6c95", x"6c97", x"6c98", x"6c9a", 
    x"6c9c", x"6c9d", x"6c9f", x"6ca1", x"6ca2", x"6ca4", x"6ca6", x"6ca7", 
    x"6ca9", x"6cab", x"6cac", x"6cae", x"6cb0", x"6cb1", x"6cb3", x"6cb5", 
    x"6cb6", x"6cb8", x"6cba", x"6cbb", x"6cbd", x"6cbf", x"6cc0", x"6cc2", 
    x"6cc3", x"6cc5", x"6cc7", x"6cc8", x"6cca", x"6ccc", x"6ccd", x"6ccf", 
    x"6cd1", x"6cd2", x"6cd4", x"6cd6", x"6cd7", x"6cd9", x"6cdb", x"6cdc", 
    x"6cde", x"6ce0", x"6ce1", x"6ce3", x"6ce5", x"6ce6", x"6ce8", x"6cea", 
    x"6ceb", x"6ced", x"6cee", x"6cf0", x"6cf2", x"6cf3", x"6cf5", x"6cf7", 
    x"6cf8", x"6cfa", x"6cfc", x"6cfd", x"6cff", x"6d01", x"6d02", x"6d04", 
    x"6d06", x"6d07", x"6d09", x"6d0a", x"6d0c", x"6d0e", x"6d0f", x"6d11", 
    x"6d13", x"6d14", x"6d16", x"6d18", x"6d19", x"6d1b", x"6d1d", x"6d1e", 
    x"6d20", x"6d21", x"6d23", x"6d25", x"6d26", x"6d28", x"6d2a", x"6d2b", 
    x"6d2d", x"6d2f", x"6d30", x"6d32", x"6d34", x"6d35", x"6d37", x"6d38", 
    x"6d3a", x"6d3c", x"6d3d", x"6d3f", x"6d41", x"6d42", x"6d44", x"6d46", 
    x"6d47", x"6d49", x"6d4a", x"6d4c", x"6d4e", x"6d4f", x"6d51", x"6d53", 
    x"6d54", x"6d56", x"6d58", x"6d59", x"6d5b", x"6d5c", x"6d5e", x"6d60", 
    x"6d61", x"6d63", x"6d65", x"6d66", x"6d68", x"6d69", x"6d6b", x"6d6d", 
    x"6d6e", x"6d70", x"6d72", x"6d73", x"6d75", x"6d76", x"6d78", x"6d7a", 
    x"6d7b", x"6d7d", x"6d7f", x"6d80", x"6d82", x"6d84", x"6d85", x"6d87", 
    x"6d88", x"6d8a", x"6d8c", x"6d8d", x"6d8f", x"6d91", x"6d92", x"6d94", 
    x"6d95", x"6d97", x"6d99", x"6d9a", x"6d9c", x"6d9d", x"6d9f", x"6da1", 
    x"6da2", x"6da4", x"6da6", x"6da7", x"6da9", x"6daa", x"6dac", x"6dae", 
    x"6daf", x"6db1", x"6db3", x"6db4", x"6db6", x"6db7", x"6db9", x"6dbb", 
    x"6dbc", x"6dbe", x"6dbf", x"6dc1", x"6dc3", x"6dc4", x"6dc6", x"6dc8", 
    x"6dc9", x"6dcb", x"6dcc", x"6dce", x"6dd0", x"6dd1", x"6dd3", x"6dd4", 
    x"6dd6", x"6dd8", x"6dd9", x"6ddb", x"6ddd", x"6dde", x"6de0", x"6de1", 
    x"6de3", x"6de5", x"6de6", x"6de8", x"6de9", x"6deb", x"6ded", x"6dee", 
    x"6df0", x"6df1", x"6df3", x"6df5", x"6df6", x"6df8", x"6dfa", x"6dfb", 
    x"6dfd", x"6dfe", x"6e00", x"6e02", x"6e03", x"6e05", x"6e06", x"6e08", 
    x"6e0a", x"6e0b", x"6e0d", x"6e0e", x"6e10", x"6e12", x"6e13", x"6e15", 
    x"6e16", x"6e18", x"6e1a", x"6e1b", x"6e1d", x"6e1e", x"6e20", x"6e22", 
    x"6e23", x"6e25", x"6e26", x"6e28", x"6e2a", x"6e2b", x"6e2d", x"6e2e", 
    x"6e30", x"6e32", x"6e33", x"6e35", x"6e36", x"6e38", x"6e3a", x"6e3b", 
    x"6e3d", x"6e3e", x"6e40", x"6e42", x"6e43", x"6e45", x"6e46", x"6e48", 
    x"6e4a", x"6e4b", x"6e4d", x"6e4e", x"6e50", x"6e52", x"6e53", x"6e55", 
    x"6e56", x"6e58", x"6e59", x"6e5b", x"6e5d", x"6e5e", x"6e60", x"6e61", 
    x"6e63", x"6e65", x"6e66", x"6e68", x"6e69", x"6e6b", x"6e6d", x"6e6e", 
    x"6e70", x"6e71", x"6e73", x"6e75", x"6e76", x"6e78", x"6e79", x"6e7b", 
    x"6e7c", x"6e7e", x"6e80", x"6e81", x"6e83", x"6e84", x"6e86", x"6e88", 
    x"6e89", x"6e8b", x"6e8c", x"6e8e", x"6e8f", x"6e91", x"6e93", x"6e94", 
    x"6e96", x"6e97", x"6e99", x"6e9b", x"6e9c", x"6e9e", x"6e9f", x"6ea1", 
    x"6ea2", x"6ea4", x"6ea6", x"6ea7", x"6ea9", x"6eaa", x"6eac", x"6ead", 
    x"6eaf", x"6eb1", x"6eb2", x"6eb4", x"6eb5", x"6eb7", x"6eb9", x"6eba", 
    x"6ebc", x"6ebd", x"6ebf", x"6ec0", x"6ec2", x"6ec4", x"6ec5", x"6ec7", 
    x"6ec8", x"6eca", x"6ecb", x"6ecd", x"6ecf", x"6ed0", x"6ed2", x"6ed3", 
    x"6ed5", x"6ed6", x"6ed8", x"6eda", x"6edb", x"6edd", x"6ede", x"6ee0", 
    x"6ee1", x"6ee3", x"6ee5", x"6ee6", x"6ee8", x"6ee9", x"6eeb", x"6eec", 
    x"6eee", x"6ef0", x"6ef1", x"6ef3", x"6ef4", x"6ef6", x"6ef7", x"6ef9", 
    x"6efb", x"6efc", x"6efe", x"6eff", x"6f01", x"6f02", x"6f04", x"6f05", 
    x"6f07", x"6f09", x"6f0a", x"6f0c", x"6f0d", x"6f0f", x"6f10", x"6f12", 
    x"6f14", x"6f15", x"6f17", x"6f18", x"6f1a", x"6f1b", x"6f1d", x"6f1e", 
    x"6f20", x"6f22", x"6f23", x"6f25", x"6f26", x"6f28", x"6f29", x"6f2b", 
    x"6f2c", x"6f2e", x"6f30", x"6f31", x"6f33", x"6f34", x"6f36", x"6f37", 
    x"6f39", x"6f3a", x"6f3c", x"6f3e", x"6f3f", x"6f41", x"6f42", x"6f44", 
    x"6f45", x"6f47", x"6f48", x"6f4a", x"6f4c", x"6f4d", x"6f4f", x"6f50", 
    x"6f52", x"6f53", x"6f55", x"6f56", x"6f58", x"6f59", x"6f5b", x"6f5d", 
    x"6f5e", x"6f60", x"6f61", x"6f63", x"6f64", x"6f66", x"6f67", x"6f69", 
    x"6f6b", x"6f6c", x"6f6e", x"6f6f", x"6f71", x"6f72", x"6f74", x"6f75", 
    x"6f77", x"6f78", x"6f7a", x"6f7c", x"6f7d", x"6f7f", x"6f80", x"6f82", 
    x"6f83", x"6f85", x"6f86", x"6f88", x"6f89", x"6f8b", x"6f8c", x"6f8e", 
    x"6f90", x"6f91", x"6f93", x"6f94", x"6f96", x"6f97", x"6f99", x"6f9a", 
    x"6f9c", x"6f9d", x"6f9f", x"6fa0", x"6fa2", x"6fa4", x"6fa5", x"6fa7", 
    x"6fa8", x"6faa", x"6fab", x"6fad", x"6fae", x"6fb0", x"6fb1", x"6fb3", 
    x"6fb4", x"6fb6", x"6fb8", x"6fb9", x"6fbb", x"6fbc", x"6fbe", x"6fbf", 
    x"6fc1", x"6fc2", x"6fc4", x"6fc5", x"6fc7", x"6fc8", x"6fca", x"6fcb", 
    x"6fcd", x"6fce", x"6fd0", x"6fd2", x"6fd3", x"6fd5", x"6fd6", x"6fd8", 
    x"6fd9", x"6fdb", x"6fdc", x"6fde", x"6fdf", x"6fe1", x"6fe2", x"6fe4", 
    x"6fe5", x"6fe7", x"6fe8", x"6fea", x"6feb", x"6fed", x"6fef", x"6ff0", 
    x"6ff2", x"6ff3", x"6ff5", x"6ff6", x"6ff8", x"6ff9", x"6ffb", x"6ffc", 
    x"6ffe", x"6fff", x"7001", x"7002", x"7004", x"7005", x"7007", x"7008", 
    x"700a", x"700b", x"700d", x"700e", x"7010", x"7012", x"7013", x"7015", 
    x"7016", x"7018", x"7019", x"701b", x"701c", x"701e", x"701f", x"7021", 
    x"7022", x"7024", x"7025", x"7027", x"7028", x"702a", x"702b", x"702d", 
    x"702e", x"7030", x"7031", x"7033", x"7034", x"7036", x"7037", x"7039", 
    x"703a", x"703c", x"703d", x"703f", x"7040", x"7042", x"7043", x"7045", 
    x"7046", x"7048", x"7049", x"704b", x"704c", x"704e", x"7050", x"7051", 
    x"7053", x"7054", x"7056", x"7057", x"7059", x"705a", x"705c", x"705d", 
    x"705f", x"7060", x"7062", x"7063", x"7065", x"7066", x"7068", x"7069", 
    x"706b", x"706c", x"706e", x"706f", x"7071", x"7072", x"7074", x"7075", 
    x"7077", x"7078", x"707a", x"707b", x"707d", x"707e", x"7080", x"7081", 
    x"7083", x"7084", x"7086", x"7087", x"7089", x"708a", x"708c", x"708d", 
    x"708f", x"7090", x"7092", x"7093", x"7095", x"7096", x"7098", x"7099", 
    x"709b", x"709c", x"709e", x"709f", x"70a0", x"70a2", x"70a3", x"70a5", 
    x"70a6", x"70a8", x"70a9", x"70ab", x"70ac", x"70ae", x"70af", x"70b1", 
    x"70b2", x"70b4", x"70b5", x"70b7", x"70b8", x"70ba", x"70bb", x"70bd", 
    x"70be", x"70c0", x"70c1", x"70c3", x"70c4", x"70c6", x"70c7", x"70c9", 
    x"70ca", x"70cc", x"70cd", x"70cf", x"70d0", x"70d2", x"70d3", x"70d5", 
    x"70d6", x"70d8", x"70d9", x"70db", x"70dc", x"70dd", x"70df", x"70e0", 
    x"70e2", x"70e3", x"70e5", x"70e6", x"70e8", x"70e9", x"70eb", x"70ec", 
    x"70ee", x"70ef", x"70f1", x"70f2", x"70f4", x"70f5", x"70f7", x"70f8", 
    x"70fa", x"70fb", x"70fd", x"70fe", x"70ff", x"7101", x"7102", x"7104", 
    x"7105", x"7107", x"7108", x"710a", x"710b", x"710d", x"710e", x"7110", 
    x"7111", x"7113", x"7114", x"7116", x"7117", x"7119", x"711a", x"711b", 
    x"711d", x"711e", x"7120", x"7121", x"7123", x"7124", x"7126", x"7127", 
    x"7129", x"712a", x"712c", x"712d", x"712f", x"7130", x"7131", x"7133", 
    x"7134", x"7136", x"7137", x"7139", x"713a", x"713c", x"713d", x"713f", 
    x"7140", x"7142", x"7143", x"7145", x"7146", x"7147", x"7149", x"714a", 
    x"714c", x"714d", x"714f", x"7150", x"7152", x"7153", x"7155", x"7156", 
    x"7158", x"7159", x"715a", x"715c", x"715d", x"715f", x"7160", x"7162", 
    x"7163", x"7165", x"7166", x"7168", x"7169", x"716a", x"716c", x"716d", 
    x"716f", x"7170", x"7172", x"7173", x"7175", x"7176", x"7178", x"7179", 
    x"717a", x"717c", x"717d", x"717f", x"7180", x"7182", x"7183", x"7185", 
    x"7186", x"7188", x"7189", x"718a", x"718c", x"718d", x"718f", x"7190", 
    x"7192", x"7193", x"7195", x"7196", x"7197", x"7199", x"719a", x"719c", 
    x"719d", x"719f", x"71a0", x"71a2", x"71a3", x"71a5", x"71a6", x"71a7", 
    x"71a9", x"71aa", x"71ac", x"71ad", x"71af", x"71b0", x"71b2", x"71b3", 
    x"71b4", x"71b6", x"71b7", x"71b9", x"71ba", x"71bc", x"71bd", x"71be", 
    x"71c0", x"71c1", x"71c3", x"71c4", x"71c6", x"71c7", x"71c9", x"71ca", 
    x"71cb", x"71cd", x"71ce", x"71d0", x"71d1", x"71d3", x"71d4", x"71d6", 
    x"71d7", x"71d8", x"71da", x"71db", x"71dd", x"71de", x"71e0", x"71e1", 
    x"71e2", x"71e4", x"71e5", x"71e7", x"71e8", x"71ea", x"71eb", x"71ec", 
    x"71ee", x"71ef", x"71f1", x"71f2", x"71f4", x"71f5", x"71f6", x"71f8", 
    x"71f9", x"71fb", x"71fc", x"71fe", x"71ff", x"7200", x"7202", x"7203", 
    x"7205", x"7206", x"7208", x"7209", x"720a", x"720c", x"720d", x"720f", 
    x"7210", x"7212", x"7213", x"7214", x"7216", x"7217", x"7219", x"721a", 
    x"721c", x"721d", x"721e", x"7220", x"7221", x"7223", x"7224", x"7226", 
    x"7227", x"7228", x"722a", x"722b", x"722d", x"722e", x"722f", x"7231", 
    x"7232", x"7234", x"7235", x"7237", x"7238", x"7239", x"723b", x"723c", 
    x"723e", x"723f", x"7240", x"7242", x"7243", x"7245", x"7246", x"7248", 
    x"7249", x"724a", x"724c", x"724d", x"724f", x"7250", x"7251", x"7253", 
    x"7254", x"7256", x"7257", x"7259", x"725a", x"725b", x"725d", x"725e", 
    x"7260", x"7261", x"7262", x"7264", x"7265", x"7267", x"7268", x"7269", 
    x"726b", x"726c", x"726e", x"726f", x"7270", x"7272", x"7273", x"7275", 
    x"7276", x"7278", x"7279", x"727a", x"727c", x"727d", x"727f", x"7280", 
    x"7281", x"7283", x"7284", x"7286", x"7287", x"7288", x"728a", x"728b", 
    x"728d", x"728e", x"728f", x"7291", x"7292", x"7294", x"7295", x"7296", 
    x"7298", x"7299", x"729b", x"729c", x"729d", x"729f", x"72a0", x"72a2", 
    x"72a3", x"72a4", x"72a6", x"72a7", x"72a9", x"72aa", x"72ab", x"72ad", 
    x"72ae", x"72b0", x"72b1", x"72b2", x"72b4", x"72b5", x"72b6", x"72b8", 
    x"72b9", x"72bb", x"72bc", x"72bd", x"72bf", x"72c0", x"72c2", x"72c3", 
    x"72c4", x"72c6", x"72c7", x"72c9", x"72ca", x"72cb", x"72cd", x"72ce", 
    x"72d0", x"72d1", x"72d2", x"72d4", x"72d5", x"72d6", x"72d8", x"72d9", 
    x"72db", x"72dc", x"72dd", x"72df", x"72e0", x"72e2", x"72e3", x"72e4", 
    x"72e6", x"72e7", x"72e8", x"72ea", x"72eb", x"72ed", x"72ee", x"72ef", 
    x"72f1", x"72f2", x"72f4", x"72f5", x"72f6", x"72f8", x"72f9", x"72fa", 
    x"72fc", x"72fd", x"72ff", x"7300", x"7301", x"7303", x"7304", x"7305", 
    x"7307", x"7308", x"730a", x"730b", x"730c", x"730e", x"730f", x"7311", 
    x"7312", x"7313", x"7315", x"7316", x"7317", x"7319", x"731a", x"731c", 
    x"731d", x"731e", x"7320", x"7321", x"7322", x"7324", x"7325", x"7326", 
    x"7328", x"7329", x"732b", x"732c", x"732d", x"732f", x"7330", x"7331", 
    x"7333", x"7334", x"7336", x"7337", x"7338", x"733a", x"733b", x"733c", 
    x"733e", x"733f", x"7340", x"7342", x"7343", x"7345", x"7346", x"7347", 
    x"7349", x"734a", x"734b", x"734d", x"734e", x"7350", x"7351", x"7352", 
    x"7354", x"7355", x"7356", x"7358", x"7359", x"735a", x"735c", x"735d", 
    x"735e", x"7360", x"7361", x"7363", x"7364", x"7365", x"7367", x"7368", 
    x"7369", x"736b", x"736c", x"736d", x"736f", x"7370", x"7372", x"7373", 
    x"7374", x"7376", x"7377", x"7378", x"737a", x"737b", x"737c", x"737e", 
    x"737f", x"7380", x"7382", x"7383", x"7384", x"7386", x"7387", x"7389", 
    x"738a", x"738b", x"738d", x"738e", x"738f", x"7391", x"7392", x"7393", 
    x"7395", x"7396", x"7397", x"7399", x"739a", x"739b", x"739d", x"739e", 
    x"739f", x"73a1", x"73a2", x"73a4", x"73a5", x"73a6", x"73a8", x"73a9", 
    x"73aa", x"73ac", x"73ad", x"73ae", x"73b0", x"73b1", x"73b2", x"73b4", 
    x"73b5", x"73b6", x"73b8", x"73b9", x"73ba", x"73bc", x"73bd", x"73be", 
    x"73c0", x"73c1", x"73c2", x"73c4", x"73c5", x"73c6", x"73c8", x"73c9", 
    x"73ca", x"73cc", x"73cd", x"73ce", x"73d0", x"73d1", x"73d3", x"73d4", 
    x"73d5", x"73d7", x"73d8", x"73d9", x"73db", x"73dc", x"73dd", x"73df", 
    x"73e0", x"73e1", x"73e3", x"73e4", x"73e5", x"73e7", x"73e8", x"73e9", 
    x"73eb", x"73ec", x"73ed", x"73ef", x"73f0", x"73f1", x"73f3", x"73f4", 
    x"73f5", x"73f7", x"73f8", x"73f9", x"73fa", x"73fc", x"73fd", x"73fe", 
    x"7400", x"7401", x"7402", x"7404", x"7405", x"7406", x"7408", x"7409", 
    x"740a", x"740c", x"740d", x"740e", x"7410", x"7411", x"7412", x"7414", 
    x"7415", x"7416", x"7418", x"7419", x"741a", x"741c", x"741d", x"741e", 
    x"7420", x"7421", x"7422", x"7424", x"7425", x"7426", x"7428", x"7429", 
    x"742a", x"742b", x"742d", x"742e", x"742f", x"7431", x"7432", x"7433", 
    x"7435", x"7436", x"7437", x"7439", x"743a", x"743b", x"743d", x"743e", 
    x"743f", x"7441", x"7442", x"7443", x"7444", x"7446", x"7447", x"7448", 
    x"744a", x"744b", x"744c", x"744e", x"744f", x"7450", x"7452", x"7453", 
    x"7454", x"7456", x"7457", x"7458", x"7459", x"745b", x"745c", x"745d", 
    x"745f", x"7460", x"7461", x"7463", x"7464", x"7465", x"7467", x"7468", 
    x"7469", x"746a", x"746c", x"746d", x"746e", x"7470", x"7471", x"7472", 
    x"7474", x"7475", x"7476", x"7478", x"7479", x"747a", x"747b", x"747d", 
    x"747e", x"747f", x"7481", x"7482", x"7483", x"7485", x"7486", x"7487", 
    x"7488", x"748a", x"748b", x"748c", x"748e", x"748f", x"7490", x"7492", 
    x"7493", x"7494", x"7495", x"7497", x"7498", x"7499", x"749b", x"749c", 
    x"749d", x"749e", x"74a0", x"74a1", x"74a2", x"74a4", x"74a5", x"74a6", 
    x"74a8", x"74a9", x"74aa", x"74ab", x"74ad", x"74ae", x"74af", x"74b1", 
    x"74b2", x"74b3", x"74b4", x"74b6", x"74b7", x"74b8", x"74ba", x"74bb", 
    x"74bc", x"74bd", x"74bf", x"74c0", x"74c1", x"74c3", x"74c4", x"74c5", 
    x"74c6", x"74c8", x"74c9", x"74ca", x"74cc", x"74cd", x"74ce", x"74cf", 
    x"74d1", x"74d2", x"74d3", x"74d5", x"74d6", x"74d7", x"74d8", x"74da", 
    x"74db", x"74dc", x"74de", x"74df", x"74e0", x"74e1", x"74e3", x"74e4", 
    x"74e5", x"74e7", x"74e8", x"74e9", x"74ea", x"74ec", x"74ed", x"74ee", 
    x"74f0", x"74f1", x"74f2", x"74f3", x"74f5", x"74f6", x"74f7", x"74f8", 
    x"74fa", x"74fb", x"74fc", x"74fe", x"74ff", x"7500", x"7501", x"7503", 
    x"7504", x"7505", x"7506", x"7508", x"7509", x"750a", x"750c", x"750d", 
    x"750e", x"750f", x"7511", x"7512", x"7513", x"7514", x"7516", x"7517", 
    x"7518", x"751a", x"751b", x"751c", x"751d", x"751f", x"7520", x"7521", 
    x"7522", x"7524", x"7525", x"7526", x"7527", x"7529", x"752a", x"752b", 
    x"752d", x"752e", x"752f", x"7530", x"7532", x"7533", x"7534", x"7535", 
    x"7537", x"7538", x"7539", x"753a", x"753c", x"753d", x"753e", x"753f", 
    x"7541", x"7542", x"7543", x"7544", x"7546", x"7547", x"7548", x"754a", 
    x"754b", x"754c", x"754d", x"754f", x"7550", x"7551", x"7552", x"7554", 
    x"7555", x"7556", x"7557", x"7559", x"755a", x"755b", x"755c", x"755e", 
    x"755f", x"7560", x"7561", x"7563", x"7564", x"7565", x"7566", x"7568", 
    x"7569", x"756a", x"756b", x"756d", x"756e", x"756f", x"7570", x"7572", 
    x"7573", x"7574", x"7575", x"7577", x"7578", x"7579", x"757a", x"757c", 
    x"757d", x"757e", x"757f", x"7581", x"7582", x"7583", x"7584", x"7586", 
    x"7587", x"7588", x"7589", x"758b", x"758c", x"758d", x"758e", x"7590", 
    x"7591", x"7592", x"7593", x"7594", x"7596", x"7597", x"7598", x"7599", 
    x"759b", x"759c", x"759d", x"759e", x"75a0", x"75a1", x"75a2", x"75a3", 
    x"75a5", x"75a6", x"75a7", x"75a8", x"75aa", x"75ab", x"75ac", x"75ad", 
    x"75ae", x"75b0", x"75b1", x"75b2", x"75b3", x"75b5", x"75b6", x"75b7", 
    x"75b8", x"75ba", x"75bb", x"75bc", x"75bd", x"75bf", x"75c0", x"75c1", 
    x"75c2", x"75c3", x"75c5", x"75c6", x"75c7", x"75c8", x"75ca", x"75cb", 
    x"75cc", x"75cd", x"75cf", x"75d0", x"75d1", x"75d2", x"75d3", x"75d5", 
    x"75d6", x"75d7", x"75d8", x"75da", x"75db", x"75dc", x"75dd", x"75de", 
    x"75e0", x"75e1", x"75e2", x"75e3", x"75e5", x"75e6", x"75e7", x"75e8", 
    x"75e9", x"75eb", x"75ec", x"75ed", x"75ee", x"75f0", x"75f1", x"75f2", 
    x"75f3", x"75f4", x"75f6", x"75f7", x"75f8", x"75f9", x"75fb", x"75fc", 
    x"75fd", x"75fe", x"75ff", x"7601", x"7602", x"7603", x"7604", x"7606", 
    x"7607", x"7608", x"7609", x"760a", x"760c", x"760d", x"760e", x"760f", 
    x"7610", x"7612", x"7613", x"7614", x"7615", x"7617", x"7618", x"7619", 
    x"761a", x"761b", x"761d", x"761e", x"761f", x"7620", x"7621", x"7623", 
    x"7624", x"7625", x"7626", x"7627", x"7629", x"762a", x"762b", x"762c", 
    x"762d", x"762f", x"7630", x"7631", x"7632", x"7634", x"7635", x"7636", 
    x"7637", x"7638", x"763a", x"763b", x"763c", x"763d", x"763e", x"7640", 
    x"7641", x"7642", x"7643", x"7644", x"7646", x"7647", x"7648", x"7649", 
    x"764a", x"764c", x"764d", x"764e", x"764f", x"7650", x"7652", x"7653", 
    x"7654", x"7655", x"7656", x"7658", x"7659", x"765a", x"765b", x"765c", 
    x"765e", x"765f", x"7660", x"7661", x"7662", x"7664", x"7665", x"7666", 
    x"7667", x"7668", x"7669", x"766b", x"766c", x"766d", x"766e", x"766f", 
    x"7671", x"7672", x"7673", x"7674", x"7675", x"7677", x"7678", x"7679", 
    x"767a", x"767b", x"767d", x"767e", x"767f", x"7680", x"7681", x"7682", 
    x"7684", x"7685", x"7686", x"7687", x"7688", x"768a", x"768b", x"768c", 
    x"768d", x"768e", x"768f", x"7691", x"7692", x"7693", x"7694", x"7695", 
    x"7697", x"7698", x"7699", x"769a", x"769b", x"769d", x"769e", x"769f", 
    x"76a0", x"76a1", x"76a2", x"76a4", x"76a5", x"76a6", x"76a7", x"76a8", 
    x"76a9", x"76ab", x"76ac", x"76ad", x"76ae", x"76af", x"76b1", x"76b2", 
    x"76b3", x"76b4", x"76b5", x"76b6", x"76b8", x"76b9", x"76ba", x"76bb", 
    x"76bc", x"76bd", x"76bf", x"76c0", x"76c1", x"76c2", x"76c3", x"76c4", 
    x"76c6", x"76c7", x"76c8", x"76c9", x"76ca", x"76cc", x"76cd", x"76ce", 
    x"76cf", x"76d0", x"76d1", x"76d3", x"76d4", x"76d5", x"76d6", x"76d7", 
    x"76d8", x"76da", x"76db", x"76dc", x"76dd", x"76de", x"76df", x"76e1", 
    x"76e2", x"76e3", x"76e4", x"76e5", x"76e6", x"76e7", x"76e9", x"76ea", 
    x"76eb", x"76ec", x"76ed", x"76ee", x"76f0", x"76f1", x"76f2", x"76f3", 
    x"76f4", x"76f5", x"76f7", x"76f8", x"76f9", x"76fa", x"76fb", x"76fc", 
    x"76fe", x"76ff", x"7700", x"7701", x"7702", x"7703", x"7704", x"7706", 
    x"7707", x"7708", x"7709", x"770a", x"770b", x"770d", x"770e", x"770f", 
    x"7710", x"7711", x"7712", x"7713", x"7715", x"7716", x"7717", x"7718", 
    x"7719", x"771a", x"771c", x"771d", x"771e", x"771f", x"7720", x"7721", 
    x"7722", x"7724", x"7725", x"7726", x"7727", x"7728", x"7729", x"772a", 
    x"772c", x"772d", x"772e", x"772f", x"7730", x"7731", x"7732", x"7734", 
    x"7735", x"7736", x"7737", x"7738", x"7739", x"773a", x"773c", x"773d", 
    x"773e", x"773f", x"7740", x"7741", x"7742", x"7744", x"7745", x"7746", 
    x"7747", x"7748", x"7749", x"774a", x"774c", x"774d", x"774e", x"774f", 
    x"7750", x"7751", x"7752", x"7754", x"7755", x"7756", x"7757", x"7758", 
    x"7759", x"775a", x"775c", x"775d", x"775e", x"775f", x"7760", x"7761", 
    x"7762", x"7763", x"7765", x"7766", x"7767", x"7768", x"7769", x"776a", 
    x"776b", x"776d", x"776e", x"776f", x"7770", x"7771", x"7772", x"7773", 
    x"7774", x"7776", x"7777", x"7778", x"7779", x"777a", x"777b", x"777c", 
    x"777d", x"777f", x"7780", x"7781", x"7782", x"7783", x"7784", x"7785", 
    x"7786", x"7788", x"7789", x"778a", x"778b", x"778c", x"778d", x"778e", 
    x"778f", x"7791", x"7792", x"7793", x"7794", x"7795", x"7796", x"7797", 
    x"7798", x"7799", x"779b", x"779c", x"779d", x"779e", x"779f", x"77a0", 
    x"77a1", x"77a2", x"77a4", x"77a5", x"77a6", x"77a7", x"77a8", x"77a9", 
    x"77aa", x"77ab", x"77ac", x"77ae", x"77af", x"77b0", x"77b1", x"77b2", 
    x"77b3", x"77b4", x"77b5", x"77b6", x"77b8", x"77b9", x"77ba", x"77bb", 
    x"77bc", x"77bd", x"77be", x"77bf", x"77c0", x"77c2", x"77c3", x"77c4", 
    x"77c5", x"77c6", x"77c7", x"77c8", x"77c9", x"77ca", x"77cc", x"77cd", 
    x"77ce", x"77cf", x"77d0", x"77d1", x"77d2", x"77d3", x"77d4", x"77d6", 
    x"77d7", x"77d8", x"77d9", x"77da", x"77db", x"77dc", x"77dd", x"77de", 
    x"77df", x"77e1", x"77e2", x"77e3", x"77e4", x"77e5", x"77e6", x"77e7", 
    x"77e8", x"77e9", x"77ea", x"77ec", x"77ed", x"77ee", x"77ef", x"77f0", 
    x"77f1", x"77f2", x"77f3", x"77f4", x"77f5", x"77f7", x"77f8", x"77f9", 
    x"77fa", x"77fb", x"77fc", x"77fd", x"77fe", x"77ff", x"7800", x"7801", 
    x"7803", x"7804", x"7805", x"7806", x"7807", x"7808", x"7809", x"780a", 
    x"780b", x"780c", x"780d", x"780f", x"7810", x"7811", x"7812", x"7813", 
    x"7814", x"7815", x"7816", x"7817", x"7818", x"7819", x"781a", x"781c", 
    x"781d", x"781e", x"781f", x"7820", x"7821", x"7822", x"7823", x"7824", 
    x"7825", x"7826", x"7828", x"7829", x"782a", x"782b", x"782c", x"782d", 
    x"782e", x"782f", x"7830", x"7831", x"7832", x"7833", x"7834", x"7836", 
    x"7837", x"7838", x"7839", x"783a", x"783b", x"783c", x"783d", x"783e", 
    x"783f", x"7840", x"7841", x"7842", x"7844", x"7845", x"7846", x"7847", 
    x"7848", x"7849", x"784a", x"784b", x"784c", x"784d", x"784e", x"784f", 
    x"7850", x"7852", x"7853", x"7854", x"7855", x"7856", x"7857", x"7858", 
    x"7859", x"785a", x"785b", x"785c", x"785d", x"785e", x"785f", x"7860", 
    x"7862", x"7863", x"7864", x"7865", x"7866", x"7867", x"7868", x"7869", 
    x"786a", x"786b", x"786c", x"786d", x"786e", x"786f", x"7870", x"7872", 
    x"7873", x"7874", x"7875", x"7876", x"7877", x"7878", x"7879", x"787a", 
    x"787b", x"787c", x"787d", x"787e", x"787f", x"7880", x"7881", x"7883", 
    x"7884", x"7885", x"7886", x"7887", x"7888", x"7889", x"788a", x"788b", 
    x"788c", x"788d", x"788e", x"788f", x"7890", x"7891", x"7892", x"7893", 
    x"7894", x"7896", x"7897", x"7898", x"7899", x"789a", x"789b", x"789c", 
    x"789d", x"789e", x"789f", x"78a0", x"78a1", x"78a2", x"78a3", x"78a4", 
    x"78a5", x"78a6", x"78a7", x"78a8", x"78a9", x"78ab", x"78ac", x"78ad", 
    x"78ae", x"78af", x"78b0", x"78b1", x"78b2", x"78b3", x"78b4", x"78b5", 
    x"78b6", x"78b7", x"78b8", x"78b9", x"78ba", x"78bb", x"78bc", x"78bd", 
    x"78be", x"78bf", x"78c0", x"78c2", x"78c3", x"78c4", x"78c5", x"78c6", 
    x"78c7", x"78c8", x"78c9", x"78ca", x"78cb", x"78cc", x"78cd", x"78ce", 
    x"78cf", x"78d0", x"78d1", x"78d2", x"78d3", x"78d4", x"78d5", x"78d6", 
    x"78d7", x"78d8", x"78d9", x"78da", x"78db", x"78dd", x"78de", x"78df", 
    x"78e0", x"78e1", x"78e2", x"78e3", x"78e4", x"78e5", x"78e6", x"78e7", 
    x"78e8", x"78e9", x"78ea", x"78eb", x"78ec", x"78ed", x"78ee", x"78ef", 
    x"78f0", x"78f1", x"78f2", x"78f3", x"78f4", x"78f5", x"78f6", x"78f7", 
    x"78f8", x"78f9", x"78fa", x"78fb", x"78fc", x"78fd", x"78fe", x"7900", 
    x"7901", x"7902", x"7903", x"7904", x"7905", x"7906", x"7907", x"7908", 
    x"7909", x"790a", x"790b", x"790c", x"790d", x"790e", x"790f", x"7910", 
    x"7911", x"7912", x"7913", x"7914", x"7915", x"7916", x"7917", x"7918", 
    x"7919", x"791a", x"791b", x"791c", x"791d", x"791e", x"791f", x"7920", 
    x"7921", x"7922", x"7923", x"7924", x"7925", x"7926", x"7927", x"7928", 
    x"7929", x"792a", x"792b", x"792c", x"792d", x"792e", x"792f", x"7930", 
    x"7931", x"7932", x"7933", x"7934", x"7935", x"7936", x"7937", x"7938", 
    x"7939", x"793a", x"793b", x"793c", x"793d", x"793e", x"793f", x"7940", 
    x"7941", x"7943", x"7944", x"7945", x"7946", x"7947", x"7948", x"7949", 
    x"794a", x"794b", x"794c", x"794d", x"794e", x"794f", x"7950", x"7951", 
    x"7952", x"7953", x"7954", x"7955", x"7956", x"7957", x"7958", x"7959", 
    x"795a", x"795b", x"795c", x"795d", x"795e", x"795f", x"7960", x"7961", 
    x"7962", x"7963", x"7964", x"7965", x"7966", x"7967", x"7968", x"7969", 
    x"796a", x"796b", x"796b", x"796c", x"796d", x"796e", x"796f", x"7970", 
    x"7971", x"7972", x"7973", x"7974", x"7975", x"7976", x"7977", x"7978", 
    x"7979", x"797a", x"797b", x"797c", x"797d", x"797e", x"797f", x"7980", 
    x"7981", x"7982", x"7983", x"7984", x"7985", x"7986", x"7987", x"7988", 
    x"7989", x"798a", x"798b", x"798c", x"798d", x"798e", x"798f", x"7990", 
    x"7991", x"7992", x"7993", x"7994", x"7995", x"7996", x"7997", x"7998", 
    x"7999", x"799a", x"799b", x"799c", x"799d", x"799e", x"799f", x"79a0", 
    x"79a1", x"79a2", x"79a3", x"79a4", x"79a5", x"79a6", x"79a7", x"79a8", 
    x"79a9", x"79aa", x"79ab", x"79ac", x"79ac", x"79ad", x"79ae", x"79af", 
    x"79b0", x"79b1", x"79b2", x"79b3", x"79b4", x"79b5", x"79b6", x"79b7", 
    x"79b8", x"79b9", x"79ba", x"79bb", x"79bc", x"79bd", x"79be", x"79bf", 
    x"79c0", x"79c1", x"79c2", x"79c3", x"79c4", x"79c5", x"79c6", x"79c7", 
    x"79c8", x"79c9", x"79ca", x"79cb", x"79cc", x"79cd", x"79cd", x"79ce", 
    x"79cf", x"79d0", x"79d1", x"79d2", x"79d3", x"79d4", x"79d5", x"79d6", 
    x"79d7", x"79d8", x"79d9", x"79da", x"79db", x"79dc", x"79dd", x"79de", 
    x"79df", x"79e0", x"79e1", x"79e2", x"79e3", x"79e4", x"79e5", x"79e6", 
    x"79e6", x"79e7", x"79e8", x"79e9", x"79ea", x"79eb", x"79ec", x"79ed", 
    x"79ee", x"79ef", x"79f0", x"79f1", x"79f2", x"79f3", x"79f4", x"79f5", 
    x"79f6", x"79f7", x"79f8", x"79f9", x"79fa", x"79fb", x"79fb", x"79fc", 
    x"79fd", x"79fe", x"79ff", x"7a00", x"7a01", x"7a02", x"7a03", x"7a04", 
    x"7a05", x"7a06", x"7a07", x"7a08", x"7a09", x"7a0a", x"7a0b", x"7a0c", 
    x"7a0d", x"7a0e", x"7a0e", x"7a0f", x"7a10", x"7a11", x"7a12", x"7a13", 
    x"7a14", x"7a15", x"7a16", x"7a17", x"7a18", x"7a19", x"7a1a", x"7a1b", 
    x"7a1c", x"7a1d", x"7a1e", x"7a1e", x"7a1f", x"7a20", x"7a21", x"7a22", 
    x"7a23", x"7a24", x"7a25", x"7a26", x"7a27", x"7a28", x"7a29", x"7a2a", 
    x"7a2b", x"7a2c", x"7a2d", x"7a2e", x"7a2e", x"7a2f", x"7a30", x"7a31", 
    x"7a32", x"7a33", x"7a34", x"7a35", x"7a36", x"7a37", x"7a38", x"7a39", 
    x"7a3a", x"7a3b", x"7a3c", x"7a3c", x"7a3d", x"7a3e", x"7a3f", x"7a40", 
    x"7a41", x"7a42", x"7a43", x"7a44", x"7a45", x"7a46", x"7a47", x"7a48", 
    x"7a49", x"7a49", x"7a4a", x"7a4b", x"7a4c", x"7a4d", x"7a4e", x"7a4f", 
    x"7a50", x"7a51", x"7a52", x"7a53", x"7a54", x"7a55", x"7a56", x"7a56", 
    x"7a57", x"7a58", x"7a59", x"7a5a", x"7a5b", x"7a5c", x"7a5d", x"7a5e", 
    x"7a5f", x"7a60", x"7a61", x"7a61", x"7a62", x"7a63", x"7a64", x"7a65", 
    x"7a66", x"7a67", x"7a68", x"7a69", x"7a6a", x"7a6b", x"7a6c", x"7a6d", 
    x"7a6d", x"7a6e", x"7a6f", x"7a70", x"7a71", x"7a72", x"7a73", x"7a74", 
    x"7a75", x"7a76", x"7a77", x"7a78", x"7a78", x"7a79", x"7a7a", x"7a7b", 
    x"7a7c", x"7a7d", x"7a7e", x"7a7f", x"7a80", x"7a81", x"7a82", x"7a82", 
    x"7a83", x"7a84", x"7a85", x"7a86", x"7a87", x"7a88", x"7a89", x"7a8a", 
    x"7a8b", x"7a8c", x"7a8c", x"7a8d", x"7a8e", x"7a8f", x"7a90", x"7a91", 
    x"7a92", x"7a93", x"7a94", x"7a95", x"7a95", x"7a96", x"7a97", x"7a98", 
    x"7a99", x"7a9a", x"7a9b", x"7a9c", x"7a9d", x"7a9e", x"7a9f", x"7a9f", 
    x"7aa0", x"7aa1", x"7aa2", x"7aa3", x"7aa4", x"7aa5", x"7aa6", x"7aa7", 
    x"7aa8", x"7aa8", x"7aa9", x"7aaa", x"7aab", x"7aac", x"7aad", x"7aae", 
    x"7aaf", x"7ab0", x"7ab0", x"7ab1", x"7ab2", x"7ab3", x"7ab4", x"7ab5", 
    x"7ab6", x"7ab7", x"7ab8", x"7ab9", x"7ab9", x"7aba", x"7abb", x"7abc", 
    x"7abd", x"7abe", x"7abf", x"7ac0", x"7ac1", x"7ac1", x"7ac2", x"7ac3", 
    x"7ac4", x"7ac5", x"7ac6", x"7ac7", x"7ac8", x"7ac9", x"7ac9", x"7aca", 
    x"7acb", x"7acc", x"7acd", x"7ace", x"7acf", x"7ad0", x"7ad1", x"7ad1", 
    x"7ad2", x"7ad3", x"7ad4", x"7ad5", x"7ad6", x"7ad7", x"7ad8", x"7ad8", 
    x"7ad9", x"7ada", x"7adb", x"7adc", x"7add", x"7ade", x"7adf", x"7ae0", 
    x"7ae0", x"7ae1", x"7ae2", x"7ae3", x"7ae4", x"7ae5", x"7ae6", x"7ae7", 
    x"7ae7", x"7ae8", x"7ae9", x"7aea", x"7aeb", x"7aec", x"7aed", x"7aee", 
    x"7aee", x"7aef", x"7af0", x"7af1", x"7af2", x"7af3", x"7af4", x"7af5", 
    x"7af5", x"7af6", x"7af7", x"7af8", x"7af9", x"7afa", x"7afb", x"7afc", 
    x"7afc", x"7afd", x"7afe", x"7aff", x"7b00", x"7b01", x"7b02", x"7b02", 
    x"7b03", x"7b04", x"7b05", x"7b06", x"7b07", x"7b08", x"7b09", x"7b09", 
    x"7b0a", x"7b0b", x"7b0c", x"7b0d", x"7b0e", x"7b0f", x"7b0f", x"7b10", 
    x"7b11", x"7b12", x"7b13", x"7b14", x"7b15", x"7b16", x"7b16", x"7b17", 
    x"7b18", x"7b19", x"7b1a", x"7b1b", x"7b1c", x"7b1c", x"7b1d", x"7b1e", 
    x"7b1f", x"7b20", x"7b21", x"7b22", x"7b22", x"7b23", x"7b24", x"7b25", 
    x"7b26", x"7b27", x"7b28", x"7b28", x"7b29", x"7b2a", x"7b2b", x"7b2c", 
    x"7b2d", x"7b2e", x"7b2e", x"7b2f", x"7b30", x"7b31", x"7b32", x"7b33", 
    x"7b33", x"7b34", x"7b35", x"7b36", x"7b37", x"7b38", x"7b39", x"7b39", 
    x"7b3a", x"7b3b", x"7b3c", x"7b3d", x"7b3e", x"7b3f", x"7b3f", x"7b40", 
    x"7b41", x"7b42", x"7b43", x"7b44", x"7b44", x"7b45", x"7b46", x"7b47", 
    x"7b48", x"7b49", x"7b4a", x"7b4a", x"7b4b", x"7b4c", x"7b4d", x"7b4e", 
    x"7b4f", x"7b4f", x"7b50", x"7b51", x"7b52", x"7b53", x"7b54", x"7b54", 
    x"7b55", x"7b56", x"7b57", x"7b58", x"7b59", x"7b5a", x"7b5a", x"7b5b", 
    x"7b5c", x"7b5d", x"7b5e", x"7b5f", x"7b5f", x"7b60", x"7b61", x"7b62", 
    x"7b63", x"7b64", x"7b64", x"7b65", x"7b66", x"7b67", x"7b68", x"7b69", 
    x"7b69", x"7b6a", x"7b6b", x"7b6c", x"7b6d", x"7b6e", x"7b6e", x"7b6f", 
    x"7b70", x"7b71", x"7b72", x"7b73", x"7b73", x"7b74", x"7b75", x"7b76", 
    x"7b77", x"7b78", x"7b78", x"7b79", x"7b7a", x"7b7b", x"7b7c", x"7b7d", 
    x"7b7d", x"7b7e", x"7b7f", x"7b80", x"7b81", x"7b81", x"7b82", x"7b83", 
    x"7b84", x"7b85", x"7b86", x"7b86", x"7b87", x"7b88", x"7b89", x"7b8a", 
    x"7b8b", x"7b8b", x"7b8c", x"7b8d", x"7b8e", x"7b8f", x"7b8f", x"7b90", 
    x"7b91", x"7b92", x"7b93", x"7b94", x"7b94", x"7b95", x"7b96", x"7b97", 
    x"7b98", x"7b98", x"7b99", x"7b9a", x"7b9b", x"7b9c", x"7b9d", x"7b9d", 
    x"7b9e", x"7b9f", x"7ba0", x"7ba1", x"7ba1", x"7ba2", x"7ba3", x"7ba4", 
    x"7ba5", x"7ba5", x"7ba6", x"7ba7", x"7ba8", x"7ba9", x"7baa", x"7baa", 
    x"7bab", x"7bac", x"7bad", x"7bae", x"7bae", x"7baf", x"7bb0", x"7bb1", 
    x"7bb2", x"7bb2", x"7bb3", x"7bb4", x"7bb5", x"7bb6", x"7bb6", x"7bb7", 
    x"7bb8", x"7bb9", x"7bba", x"7bba", x"7bbb", x"7bbc", x"7bbd", x"7bbe", 
    x"7bbf", x"7bbf", x"7bc0", x"7bc1", x"7bc2", x"7bc3", x"7bc3", x"7bc4", 
    x"7bc5", x"7bc6", x"7bc7", x"7bc7", x"7bc8", x"7bc9", x"7bca", x"7bcb", 
    x"7bcb", x"7bcc", x"7bcd", x"7bce", x"7bcf", x"7bcf", x"7bd0", x"7bd1", 
    x"7bd2", x"7bd2", x"7bd3", x"7bd4", x"7bd5", x"7bd6", x"7bd6", x"7bd7", 
    x"7bd8", x"7bd9", x"7bda", x"7bda", x"7bdb", x"7bdc", x"7bdd", x"7bde", 
    x"7bde", x"7bdf", x"7be0", x"7be1", x"7be2", x"7be2", x"7be3", x"7be4", 
    x"7be5", x"7be6", x"7be6", x"7be7", x"7be8", x"7be9", x"7be9", x"7bea", 
    x"7beb", x"7bec", x"7bed", x"7bed", x"7bee", x"7bef", x"7bf0", x"7bf1", 
    x"7bf1", x"7bf2", x"7bf3", x"7bf4", x"7bf4", x"7bf5", x"7bf6", x"7bf7", 
    x"7bf8", x"7bf8", x"7bf9", x"7bfa", x"7bfb", x"7bfb", x"7bfc", x"7bfd", 
    x"7bfe", x"7bff", x"7bff", x"7c00", x"7c01", x"7c02", x"7c02", x"7c03", 
    x"7c04", x"7c05", x"7c06", x"7c06", x"7c07", x"7c08", x"7c09", x"7c09", 
    x"7c0a", x"7c0b", x"7c0c", x"7c0d", x"7c0d", x"7c0e", x"7c0f", x"7c10", 
    x"7c10", x"7c11", x"7c12", x"7c13", x"7c14", x"7c14", x"7c15", x"7c16", 
    x"7c17", x"7c17", x"7c18", x"7c19", x"7c1a", x"7c1a", x"7c1b", x"7c1c", 
    x"7c1d", x"7c1e", x"7c1e", x"7c1f", x"7c20", x"7c21", x"7c21", x"7c22", 
    x"7c23", x"7c24", x"7c24", x"7c25", x"7c26", x"7c27", x"7c27", x"7c28", 
    x"7c29", x"7c2a", x"7c2b", x"7c2b", x"7c2c", x"7c2d", x"7c2e", x"7c2e", 
    x"7c2f", x"7c30", x"7c31", x"7c31", x"7c32", x"7c33", x"7c34", x"7c34", 
    x"7c35", x"7c36", x"7c37", x"7c37", x"7c38", x"7c39", x"7c3a", x"7c3a", 
    x"7c3b", x"7c3c", x"7c3d", x"7c3e", x"7c3e", x"7c3f", x"7c40", x"7c41", 
    x"7c41", x"7c42", x"7c43", x"7c44", x"7c44", x"7c45", x"7c46", x"7c47", 
    x"7c47", x"7c48", x"7c49", x"7c4a", x"7c4a", x"7c4b", x"7c4c", x"7c4d", 
    x"7c4d", x"7c4e", x"7c4f", x"7c50", x"7c50", x"7c51", x"7c52", x"7c53", 
    x"7c53", x"7c54", x"7c55", x"7c56", x"7c56", x"7c57", x"7c58", x"7c59", 
    x"7c59", x"7c5a", x"7c5b", x"7c5c", x"7c5c", x"7c5d", x"7c5e", x"7c5e", 
    x"7c5f", x"7c60", x"7c61", x"7c61", x"7c62", x"7c63", x"7c64", x"7c64", 
    x"7c65", x"7c66", x"7c67", x"7c67", x"7c68", x"7c69", x"7c6a", x"7c6a", 
    x"7c6b", x"7c6c", x"7c6d", x"7c6d", x"7c6e", x"7c6f", x"7c6f", x"7c70", 
    x"7c71", x"7c72", x"7c72", x"7c73", x"7c74", x"7c75", x"7c75", x"7c76", 
    x"7c77", x"7c78", x"7c78", x"7c79", x"7c7a", x"7c7a", x"7c7b", x"7c7c", 
    x"7c7d", x"7c7d", x"7c7e", x"7c7f", x"7c80", x"7c80", x"7c81", x"7c82", 
    x"7c83", x"7c83", x"7c84", x"7c85", x"7c85", x"7c86", x"7c87", x"7c88", 
    x"7c88", x"7c89", x"7c8a", x"7c8a", x"7c8b", x"7c8c", x"7c8d", x"7c8d", 
    x"7c8e", x"7c8f", x"7c90", x"7c90", x"7c91", x"7c92", x"7c92", x"7c93", 
    x"7c94", x"7c95", x"7c95", x"7c96", x"7c97", x"7c98", x"7c98", x"7c99", 
    x"7c9a", x"7c9a", x"7c9b", x"7c9c", x"7c9d", x"7c9d", x"7c9e", x"7c9f", 
    x"7c9f", x"7ca0", x"7ca1", x"7ca2", x"7ca2", x"7ca3", x"7ca4", x"7ca4", 
    x"7ca5", x"7ca6", x"7ca7", x"7ca7", x"7ca8", x"7ca9", x"7ca9", x"7caa", 
    x"7cab", x"7cac", x"7cac", x"7cad", x"7cae", x"7cae", x"7caf", x"7cb0", 
    x"7cb1", x"7cb1", x"7cb2", x"7cb3", x"7cb3", x"7cb4", x"7cb5", x"7cb5", 
    x"7cb6", x"7cb7", x"7cb8", x"7cb8", x"7cb9", x"7cba", x"7cba", x"7cbb", 
    x"7cbc", x"7cbd", x"7cbd", x"7cbe", x"7cbf", x"7cbf", x"7cc0", x"7cc1", 
    x"7cc1", x"7cc2", x"7cc3", x"7cc4", x"7cc4", x"7cc5", x"7cc6", x"7cc6", 
    x"7cc7", x"7cc8", x"7cc8", x"7cc9", x"7cca", x"7ccb", x"7ccb", x"7ccc", 
    x"7ccd", x"7ccd", x"7cce", x"7ccf", x"7ccf", x"7cd0", x"7cd1", x"7cd2", 
    x"7cd2", x"7cd3", x"7cd4", x"7cd4", x"7cd5", x"7cd6", x"7cd6", x"7cd7", 
    x"7cd8", x"7cd8", x"7cd9", x"7cda", x"7cdb", x"7cdb", x"7cdc", x"7cdd", 
    x"7cdd", x"7cde", x"7cdf", x"7cdf", x"7ce0", x"7ce1", x"7ce1", x"7ce2", 
    x"7ce3", x"7ce4", x"7ce4", x"7ce5", x"7ce6", x"7ce6", x"7ce7", x"7ce8", 
    x"7ce8", x"7ce9", x"7cea", x"7cea", x"7ceb", x"7cec", x"7cec", x"7ced", 
    x"7cee", x"7cee", x"7cef", x"7cf0", x"7cf1", x"7cf1", x"7cf2", x"7cf3", 
    x"7cf3", x"7cf4", x"7cf5", x"7cf5", x"7cf6", x"7cf7", x"7cf7", x"7cf8", 
    x"7cf9", x"7cf9", x"7cfa", x"7cfb", x"7cfb", x"7cfc", x"7cfd", x"7cfd", 
    x"7cfe", x"7cff", x"7cff", x"7d00", x"7d01", x"7d02", x"7d02", x"7d03", 
    x"7d04", x"7d04", x"7d05", x"7d06", x"7d06", x"7d07", x"7d08", x"7d08", 
    x"7d09", x"7d0a", x"7d0a", x"7d0b", x"7d0c", x"7d0c", x"7d0d", x"7d0e", 
    x"7d0e", x"7d0f", x"7d10", x"7d10", x"7d11", x"7d12", x"7d12", x"7d13", 
    x"7d14", x"7d14", x"7d15", x"7d16", x"7d16", x"7d17", x"7d18", x"7d18", 
    x"7d19", x"7d1a", x"7d1a", x"7d1b", x"7d1c", x"7d1c", x"7d1d", x"7d1e", 
    x"7d1e", x"7d1f", x"7d20", x"7d20", x"7d21", x"7d22", x"7d22", x"7d23", 
    x"7d24", x"7d24", x"7d25", x"7d26", x"7d26", x"7d27", x"7d28", x"7d28", 
    x"7d29", x"7d29", x"7d2a", x"7d2b", x"7d2b", x"7d2c", x"7d2d", x"7d2d", 
    x"7d2e", x"7d2f", x"7d2f", x"7d30", x"7d31", x"7d31", x"7d32", x"7d33", 
    x"7d33", x"7d34", x"7d35", x"7d35", x"7d36", x"7d37", x"7d37", x"7d38", 
    x"7d39", x"7d39", x"7d3a", x"7d3a", x"7d3b", x"7d3c", x"7d3c", x"7d3d", 
    x"7d3e", x"7d3e", x"7d3f", x"7d40", x"7d40", x"7d41", x"7d42", x"7d42", 
    x"7d43", x"7d44", x"7d44", x"7d45", x"7d45", x"7d46", x"7d47", x"7d47", 
    x"7d48", x"7d49", x"7d49", x"7d4a", x"7d4b", x"7d4b", x"7d4c", x"7d4d", 
    x"7d4d", x"7d4e", x"7d4e", x"7d4f", x"7d50", x"7d50", x"7d51", x"7d52", 
    x"7d52", x"7d53", x"7d54", x"7d54", x"7d55", x"7d56", x"7d56", x"7d57", 
    x"7d57", x"7d58", x"7d59", x"7d59", x"7d5a", x"7d5b", x"7d5b", x"7d5c", 
    x"7d5c", x"7d5d", x"7d5e", x"7d5e", x"7d5f", x"7d60", x"7d60", x"7d61", 
    x"7d62", x"7d62", x"7d63", x"7d63", x"7d64", x"7d65", x"7d65", x"7d66", 
    x"7d67", x"7d67", x"7d68", x"7d68", x"7d69", x"7d6a", x"7d6a", x"7d6b", 
    x"7d6c", x"7d6c", x"7d6d", x"7d6e", x"7d6e", x"7d6f", x"7d6f", x"7d70", 
    x"7d71", x"7d71", x"7d72", x"7d73", x"7d73", x"7d74", x"7d74", x"7d75", 
    x"7d76", x"7d76", x"7d77", x"7d77", x"7d78", x"7d79", x"7d79", x"7d7a", 
    x"7d7b", x"7d7b", x"7d7c", x"7d7c", x"7d7d", x"7d7e", x"7d7e", x"7d7f", 
    x"7d80", x"7d80", x"7d81", x"7d81", x"7d82", x"7d83", x"7d83", x"7d84", 
    x"7d84", x"7d85", x"7d86", x"7d86", x"7d87", x"7d88", x"7d88", x"7d89", 
    x"7d89", x"7d8a", x"7d8b", x"7d8b", x"7d8c", x"7d8c", x"7d8d", x"7d8e", 
    x"7d8e", x"7d8f", x"7d90", x"7d90", x"7d91", x"7d91", x"7d92", x"7d93", 
    x"7d93", x"7d94", x"7d94", x"7d95", x"7d96", x"7d96", x"7d97", x"7d97", 
    x"7d98", x"7d99", x"7d99", x"7d9a", x"7d9a", x"7d9b", x"7d9c", x"7d9c", 
    x"7d9d", x"7d9d", x"7d9e", x"7d9f", x"7d9f", x"7da0", x"7da0", x"7da1", 
    x"7da2", x"7da2", x"7da3", x"7da3", x"7da4", x"7da5", x"7da5", x"7da6", 
    x"7da6", x"7da7", x"7da8", x"7da8", x"7da9", x"7da9", x"7daa", x"7dab", 
    x"7dab", x"7dac", x"7dac", x"7dad", x"7dae", x"7dae", x"7daf", x"7daf", 
    x"7db0", x"7db1", x"7db1", x"7db2", x"7db2", x"7db3", x"7db4", x"7db4", 
    x"7db5", x"7db5", x"7db6", x"7db7", x"7db7", x"7db8", x"7db8", x"7db9", 
    x"7db9", x"7dba", x"7dbb", x"7dbb", x"7dbc", x"7dbc", x"7dbd", x"7dbe", 
    x"7dbe", x"7dbf", x"7dbf", x"7dc0", x"7dc1", x"7dc1", x"7dc2", x"7dc2", 
    x"7dc3", x"7dc3", x"7dc4", x"7dc5", x"7dc5", x"7dc6", x"7dc6", x"7dc7", 
    x"7dc8", x"7dc8", x"7dc9", x"7dc9", x"7dca", x"7dca", x"7dcb", x"7dcc", 
    x"7dcc", x"7dcd", x"7dcd", x"7dce", x"7dce", x"7dcf", x"7dd0", x"7dd0", 
    x"7dd1", x"7dd1", x"7dd2", x"7dd3", x"7dd3", x"7dd4", x"7dd4", x"7dd5", 
    x"7dd5", x"7dd6", x"7dd7", x"7dd7", x"7dd8", x"7dd8", x"7dd9", x"7dd9", 
    x"7dda", x"7ddb", x"7ddb", x"7ddc", x"7ddc", x"7ddd", x"7ddd", x"7dde", 
    x"7ddf", x"7ddf", x"7de0", x"7de0", x"7de1", x"7de1", x"7de2", x"7de3", 
    x"7de3", x"7de4", x"7de4", x"7de5", x"7de5", x"7de6", x"7de7", x"7de7", 
    x"7de8", x"7de8", x"7de9", x"7de9", x"7dea", x"7dea", x"7deb", x"7dec", 
    x"7dec", x"7ded", x"7ded", x"7dee", x"7dee", x"7def", x"7df0", x"7df0", 
    x"7df1", x"7df1", x"7df2", x"7df2", x"7df3", x"7df3", x"7df4", x"7df5", 
    x"7df5", x"7df6", x"7df6", x"7df7", x"7df7", x"7df8", x"7df8", x"7df9", 
    x"7dfa", x"7dfa", x"7dfb", x"7dfb", x"7dfc", x"7dfc", x"7dfd", x"7dfd", 
    x"7dfe", x"7dff", x"7dff", x"7e00", x"7e00", x"7e01", x"7e01", x"7e02", 
    x"7e02", x"7e03", x"7e04", x"7e04", x"7e05", x"7e05", x"7e06", x"7e06", 
    x"7e07", x"7e07", x"7e08", x"7e09", x"7e09", x"7e0a", x"7e0a", x"7e0b", 
    x"7e0b", x"7e0c", x"7e0c", x"7e0d", x"7e0d", x"7e0e", x"7e0f", x"7e0f", 
    x"7e10", x"7e10", x"7e11", x"7e11", x"7e12", x"7e12", x"7e13", x"7e13", 
    x"7e14", x"7e15", x"7e15", x"7e16", x"7e16", x"7e17", x"7e17", x"7e18", 
    x"7e18", x"7e19", x"7e19", x"7e1a", x"7e1a", x"7e1b", x"7e1c", x"7e1c", 
    x"7e1d", x"7e1d", x"7e1e", x"7e1e", x"7e1f", x"7e1f", x"7e20", x"7e20", 
    x"7e21", x"7e21", x"7e22", x"7e22", x"7e23", x"7e24", x"7e24", x"7e25", 
    x"7e25", x"7e26", x"7e26", x"7e27", x"7e27", x"7e28", x"7e28", x"7e29", 
    x"7e29", x"7e2a", x"7e2a", x"7e2b", x"7e2c", x"7e2c", x"7e2d", x"7e2d", 
    x"7e2e", x"7e2e", x"7e2f", x"7e2f", x"7e30", x"7e30", x"7e31", x"7e31", 
    x"7e32", x"7e32", x"7e33", x"7e33", x"7e34", x"7e34", x"7e35", x"7e36", 
    x"7e36", x"7e37", x"7e37", x"7e38", x"7e38", x"7e39", x"7e39", x"7e3a", 
    x"7e3a", x"7e3b", x"7e3b", x"7e3c", x"7e3c", x"7e3d", x"7e3d", x"7e3e", 
    x"7e3e", x"7e3f", x"7e3f", x"7e40", x"7e40", x"7e41", x"7e41", x"7e42", 
    x"7e42", x"7e43", x"7e44", x"7e44", x"7e45", x"7e45", x"7e46", x"7e46", 
    x"7e47", x"7e47", x"7e48", x"7e48", x"7e49", x"7e49", x"7e4a", x"7e4a", 
    x"7e4b", x"7e4b", x"7e4c", x"7e4c", x"7e4d", x"7e4d", x"7e4e", x"7e4e", 
    x"7e4f", x"7e4f", x"7e50", x"7e50", x"7e51", x"7e51", x"7e52", x"7e52", 
    x"7e53", x"7e53", x"7e54", x"7e54", x"7e55", x"7e55", x"7e56", x"7e56", 
    x"7e57", x"7e57", x"7e58", x"7e58", x"7e59", x"7e59", x"7e5a", x"7e5a", 
    x"7e5b", x"7e5b", x"7e5c", x"7e5c", x"7e5d", x"7e5d", x"7e5e", x"7e5e", 
    x"7e5f", x"7e5f", x"7e60", x"7e60", x"7e61", x"7e61", x"7e62", x"7e62", 
    x"7e63", x"7e63", x"7e64", x"7e64", x"7e65", x"7e65", x"7e66", x"7e66", 
    x"7e67", x"7e67", x"7e68", x"7e68", x"7e69", x"7e69", x"7e6a", x"7e6a", 
    x"7e6b", x"7e6b", x"7e6c", x"7e6c", x"7e6d", x"7e6d", x"7e6e", x"7e6e", 
    x"7e6f", x"7e6f", x"7e70", x"7e70", x"7e71", x"7e71", x"7e72", x"7e72", 
    x"7e73", x"7e73", x"7e74", x"7e74", x"7e75", x"7e75", x"7e76", x"7e76", 
    x"7e77", x"7e77", x"7e77", x"7e78", x"7e78", x"7e79", x"7e79", x"7e7a", 
    x"7e7a", x"7e7b", x"7e7b", x"7e7c", x"7e7c", x"7e7d", x"7e7d", x"7e7e", 
    x"7e7e", x"7e7f", x"7e7f", x"7e80", x"7e80", x"7e81", x"7e81", x"7e82", 
    x"7e82", x"7e83", x"7e83", x"7e83", x"7e84", x"7e84", x"7e85", x"7e85", 
    x"7e86", x"7e86", x"7e87", x"7e87", x"7e88", x"7e88", x"7e89", x"7e89", 
    x"7e8a", x"7e8a", x"7e8b", x"7e8b", x"7e8c", x"7e8c", x"7e8d", x"7e8d", 
    x"7e8d", x"7e8e", x"7e8e", x"7e8f", x"7e8f", x"7e90", x"7e90", x"7e91", 
    x"7e91", x"7e92", x"7e92", x"7e93", x"7e93", x"7e94", x"7e94", x"7e94", 
    x"7e95", x"7e95", x"7e96", x"7e96", x"7e97", x"7e97", x"7e98", x"7e98", 
    x"7e99", x"7e99", x"7e9a", x"7e9a", x"7e9b", x"7e9b", x"7e9b", x"7e9c", 
    x"7e9c", x"7e9d", x"7e9d", x"7e9e", x"7e9e", x"7e9f", x"7e9f", x"7ea0", 
    x"7ea0", x"7ea0", x"7ea1", x"7ea1", x"7ea2", x"7ea2", x"7ea3", x"7ea3", 
    x"7ea4", x"7ea4", x"7ea5", x"7ea5", x"7ea6", x"7ea6", x"7ea6", x"7ea7", 
    x"7ea7", x"7ea8", x"7ea8", x"7ea9", x"7ea9", x"7eaa", x"7eaa", x"7eaa", 
    x"7eab", x"7eab", x"7eac", x"7eac", x"7ead", x"7ead", x"7eae", x"7eae", 
    x"7eaf", x"7eaf", x"7eaf", x"7eb0", x"7eb0", x"7eb1", x"7eb1", x"7eb2", 
    x"7eb2", x"7eb3", x"7eb3", x"7eb3", x"7eb4", x"7eb4", x"7eb5", x"7eb5", 
    x"7eb6", x"7eb6", x"7eb7", x"7eb7", x"7eb7", x"7eb8", x"7eb8", x"7eb9", 
    x"7eb9", x"7eba", x"7eba", x"7ebb", x"7ebb", x"7ebb", x"7ebc", x"7ebc", 
    x"7ebd", x"7ebd", x"7ebe", x"7ebe", x"7ebf", x"7ebf", x"7ebf", x"7ec0", 
    x"7ec0", x"7ec1", x"7ec1", x"7ec2", x"7ec2", x"7ec2", x"7ec3", x"7ec3", 
    x"7ec4", x"7ec4", x"7ec5", x"7ec5", x"7ec5", x"7ec6", x"7ec6", x"7ec7", 
    x"7ec7", x"7ec8", x"7ec8", x"7ec9", x"7ec9", x"7ec9", x"7eca", x"7eca", 
    x"7ecb", x"7ecb", x"7ecc", x"7ecc", x"7ecc", x"7ecd", x"7ecd", x"7ece", 
    x"7ece", x"7ecf", x"7ecf", x"7ecf", x"7ed0", x"7ed0", x"7ed1", x"7ed1", 
    x"7ed2", x"7ed2", x"7ed2", x"7ed3", x"7ed3", x"7ed4", x"7ed4", x"7ed4", 
    x"7ed5", x"7ed5", x"7ed6", x"7ed6", x"7ed7", x"7ed7", x"7ed7", x"7ed8", 
    x"7ed8", x"7ed9", x"7ed9", x"7eda", x"7eda", x"7eda", x"7edb", x"7edb", 
    x"7edc", x"7edc", x"7edc", x"7edd", x"7edd", x"7ede", x"7ede", x"7edf", 
    x"7edf", x"7edf", x"7ee0", x"7ee0", x"7ee1", x"7ee1", x"7ee1", x"7ee2", 
    x"7ee2", x"7ee3", x"7ee3", x"7ee4", x"7ee4", x"7ee4", x"7ee5", x"7ee5", 
    x"7ee6", x"7ee6", x"7ee6", x"7ee7", x"7ee7", x"7ee8", x"7ee8", x"7ee8", 
    x"7ee9", x"7ee9", x"7eea", x"7eea", x"7eea", x"7eeb", x"7eeb", x"7eec", 
    x"7eec", x"7eed", x"7eed", x"7eed", x"7eee", x"7eee", x"7eef", x"7eef", 
    x"7eef", x"7ef0", x"7ef0", x"7ef1", x"7ef1", x"7ef1", x"7ef2", x"7ef2", 
    x"7ef3", x"7ef3", x"7ef3", x"7ef4", x"7ef4", x"7ef5", x"7ef5", x"7ef5", 
    x"7ef6", x"7ef6", x"7ef7", x"7ef7", x"7ef7", x"7ef8", x"7ef8", x"7ef9", 
    x"7ef9", x"7ef9", x"7efa", x"7efa", x"7efb", x"7efb", x"7efb", x"7efc", 
    x"7efc", x"7efd", x"7efd", x"7efd", x"7efe", x"7efe", x"7efe", x"7eff", 
    x"7eff", x"7f00", x"7f00", x"7f00", x"7f01", x"7f01", x"7f02", x"7f02", 
    x"7f02", x"7f03", x"7f03", x"7f04", x"7f04", x"7f04", x"7f05", x"7f05", 
    x"7f05", x"7f06", x"7f06", x"7f07", x"7f07", x"7f07", x"7f08", x"7f08", 
    x"7f09", x"7f09", x"7f09", x"7f0a", x"7f0a", x"7f0a", x"7f0b", x"7f0b", 
    x"7f0c", x"7f0c", x"7f0c", x"7f0d", x"7f0d", x"7f0e", x"7f0e", x"7f0e", 
    x"7f0f", x"7f0f", x"7f0f", x"7f10", x"7f10", x"7f11", x"7f11", x"7f11", 
    x"7f12", x"7f12", x"7f12", x"7f13", x"7f13", x"7f14", x"7f14", x"7f14", 
    x"7f15", x"7f15", x"7f15", x"7f16", x"7f16", x"7f17", x"7f17", x"7f17", 
    x"7f18", x"7f18", x"7f18", x"7f19", x"7f19", x"7f1a", x"7f1a", x"7f1a", 
    x"7f1b", x"7f1b", x"7f1b", x"7f1c", x"7f1c", x"7f1d", x"7f1d", x"7f1d", 
    x"7f1e", x"7f1e", x"7f1e", x"7f1f", x"7f1f", x"7f1f", x"7f20", x"7f20", 
    x"7f21", x"7f21", x"7f21", x"7f22", x"7f22", x"7f22", x"7f23", x"7f23", 
    x"7f23", x"7f24", x"7f24", x"7f25", x"7f25", x"7f25", x"7f26", x"7f26", 
    x"7f26", x"7f27", x"7f27", x"7f27", x"7f28", x"7f28", x"7f29", x"7f29", 
    x"7f29", x"7f2a", x"7f2a", x"7f2a", x"7f2b", x"7f2b", x"7f2b", x"7f2c", 
    x"7f2c", x"7f2c", x"7f2d", x"7f2d", x"7f2e", x"7f2e", x"7f2e", x"7f2f", 
    x"7f2f", x"7f2f", x"7f30", x"7f30", x"7f30", x"7f31", x"7f31", x"7f31", 
    x"7f32", x"7f32", x"7f32", x"7f33", x"7f33", x"7f34", x"7f34", x"7f34", 
    x"7f35", x"7f35", x"7f35", x"7f36", x"7f36", x"7f36", x"7f37", x"7f37", 
    x"7f37", x"7f38", x"7f38", x"7f38", x"7f39", x"7f39", x"7f39", x"7f3a", 
    x"7f3a", x"7f3a", x"7f3b", x"7f3b", x"7f3b", x"7f3c", x"7f3c", x"7f3d", 
    x"7f3d", x"7f3d", x"7f3e", x"7f3e", x"7f3e", x"7f3f", x"7f3f", x"7f3f", 
    x"7f40", x"7f40", x"7f40", x"7f41", x"7f41", x"7f41", x"7f42", x"7f42", 
    x"7f42", x"7f43", x"7f43", x"7f43", x"7f44", x"7f44", x"7f44", x"7f45", 
    x"7f45", x"7f45", x"7f46", x"7f46", x"7f46", x"7f47", x"7f47", x"7f47", 
    x"7f48", x"7f48", x"7f48", x"7f49", x"7f49", x"7f49", x"7f4a", x"7f4a", 
    x"7f4a", x"7f4b", x"7f4b", x"7f4b", x"7f4c", x"7f4c", x"7f4c", x"7f4d", 
    x"7f4d", x"7f4d", x"7f4e", x"7f4e", x"7f4e", x"7f4f", x"7f4f", x"7f4f", 
    x"7f50", x"7f50", x"7f50", x"7f50", x"7f51", x"7f51", x"7f51", x"7f52", 
    x"7f52", x"7f52", x"7f53", x"7f53", x"7f53", x"7f54", x"7f54", x"7f54", 
    x"7f55", x"7f55", x"7f55", x"7f56", x"7f56", x"7f56", x"7f57", x"7f57", 
    x"7f57", x"7f58", x"7f58", x"7f58", x"7f58", x"7f59", x"7f59", x"7f59", 
    x"7f5a", x"7f5a", x"7f5a", x"7f5b", x"7f5b", x"7f5b", x"7f5c", x"7f5c", 
    x"7f5c", x"7f5d", x"7f5d", x"7f5d", x"7f5e", x"7f5e", x"7f5e", x"7f5e", 
    x"7f5f", x"7f5f", x"7f5f", x"7f60", x"7f60", x"7f60", x"7f61", x"7f61", 
    x"7f61", x"7f62", x"7f62", x"7f62", x"7f62", x"7f63", x"7f63", x"7f63", 
    x"7f64", x"7f64", x"7f64", x"7f65", x"7f65", x"7f65", x"7f65", x"7f66", 
    x"7f66", x"7f66", x"7f67", x"7f67", x"7f67", x"7f68", x"7f68", x"7f68", 
    x"7f69", x"7f69", x"7f69", x"7f69", x"7f6a", x"7f6a", x"7f6a", x"7f6b", 
    x"7f6b", x"7f6b", x"7f6c", x"7f6c", x"7f6c", x"7f6c", x"7f6d", x"7f6d", 
    x"7f6d", x"7f6e", x"7f6e", x"7f6e", x"7f6e", x"7f6f", x"7f6f", x"7f6f", 
    x"7f70", x"7f70", x"7f70", x"7f71", x"7f71", x"7f71", x"7f71", x"7f72", 
    x"7f72", x"7f72", x"7f73", x"7f73", x"7f73", x"7f73", x"7f74", x"7f74", 
    x"7f74", x"7f75", x"7f75", x"7f75", x"7f75", x"7f76", x"7f76", x"7f76", 
    x"7f77", x"7f77", x"7f77", x"7f77", x"7f78", x"7f78", x"7f78", x"7f79", 
    x"7f79", x"7f79", x"7f79", x"7f7a", x"7f7a", x"7f7a", x"7f7b", x"7f7b", 
    x"7f7b", x"7f7b", x"7f7c", x"7f7c", x"7f7c", x"7f7d", x"7f7d", x"7f7d", 
    x"7f7d", x"7f7e", x"7f7e", x"7f7e", x"7f7f", x"7f7f", x"7f7f", x"7f7f", 
    x"7f80", x"7f80", x"7f80", x"7f80", x"7f81", x"7f81", x"7f81", x"7f82", 
    x"7f82", x"7f82", x"7f82", x"7f83", x"7f83", x"7f83", x"7f83", x"7f84", 
    x"7f84", x"7f84", x"7f85", x"7f85", x"7f85", x"7f85", x"7f86", x"7f86", 
    x"7f86", x"7f86", x"7f87", x"7f87", x"7f87", x"7f88", x"7f88", x"7f88", 
    x"7f88", x"7f89", x"7f89", x"7f89", x"7f89", x"7f8a", x"7f8a", x"7f8a", 
    x"7f8a", x"7f8b", x"7f8b", x"7f8b", x"7f8c", x"7f8c", x"7f8c", x"7f8c", 
    x"7f8d", x"7f8d", x"7f8d", x"7f8d", x"7f8e", x"7f8e", x"7f8e", x"7f8e", 
    x"7f8f", x"7f8f", x"7f8f", x"7f8f", x"7f90", x"7f90", x"7f90", x"7f90", 
    x"7f91", x"7f91", x"7f91", x"7f91", x"7f92", x"7f92", x"7f92", x"7f93", 
    x"7f93", x"7f93", x"7f93", x"7f94", x"7f94", x"7f94", x"7f94", x"7f95", 
    x"7f95", x"7f95", x"7f95", x"7f96", x"7f96", x"7f96", x"7f96", x"7f97", 
    x"7f97", x"7f97", x"7f97", x"7f98", x"7f98", x"7f98", x"7f98", x"7f99", 
    x"7f99", x"7f99", x"7f99", x"7f9a", x"7f9a", x"7f9a", x"7f9a", x"7f9b", 
    x"7f9b", x"7f9b", x"7f9b", x"7f9c", x"7f9c", x"7f9c", x"7f9c", x"7f9c", 
    x"7f9d", x"7f9d", x"7f9d", x"7f9d", x"7f9e", x"7f9e", x"7f9e", x"7f9e", 
    x"7f9f", x"7f9f", x"7f9f", x"7f9f", x"7fa0", x"7fa0", x"7fa0", x"7fa0", 
    x"7fa1", x"7fa1", x"7fa1", x"7fa1", x"7fa2", x"7fa2", x"7fa2", x"7fa2", 
    x"7fa2", x"7fa3", x"7fa3", x"7fa3", x"7fa3", x"7fa4", x"7fa4", x"7fa4", 
    x"7fa4", x"7fa5", x"7fa5", x"7fa5", x"7fa5", x"7fa6", x"7fa6", x"7fa6", 
    x"7fa6", x"7fa6", x"7fa7", x"7fa7", x"7fa7", x"7fa7", x"7fa8", x"7fa8", 
    x"7fa8", x"7fa8", x"7fa9", x"7fa9", x"7fa9", x"7fa9", x"7fa9", x"7faa", 
    x"7faa", x"7faa", x"7faa", x"7fab", x"7fab", x"7fab", x"7fab", x"7fab", 
    x"7fac", x"7fac", x"7fac", x"7fac", x"7fad", x"7fad", x"7fad", x"7fad", 
    x"7fad", x"7fae", x"7fae", x"7fae", x"7fae", x"7faf", x"7faf", x"7faf", 
    x"7faf", x"7faf", x"7fb0", x"7fb0", x"7fb0", x"7fb0", x"7fb1", x"7fb1", 
    x"7fb1", x"7fb1", x"7fb1", x"7fb2", x"7fb2", x"7fb2", x"7fb2", x"7fb2", 
    x"7fb3", x"7fb3", x"7fb3", x"7fb3", x"7fb4", x"7fb4", x"7fb4", x"7fb4", 
    x"7fb4", x"7fb5", x"7fb5", x"7fb5", x"7fb5", x"7fb5", x"7fb6", x"7fb6", 
    x"7fb6", x"7fb6", x"7fb6", x"7fb7", x"7fb7", x"7fb7", x"7fb7", x"7fb8", 
    x"7fb8", x"7fb8", x"7fb8", x"7fb8", x"7fb9", x"7fb9", x"7fb9", x"7fb9", 
    x"7fb9", x"7fba", x"7fba", x"7fba", x"7fba", x"7fba", x"7fbb", x"7fbb", 
    x"7fbb", x"7fbb", x"7fbb", x"7fbc", x"7fbc", x"7fbc", x"7fbc", x"7fbc", 
    x"7fbd", x"7fbd", x"7fbd", x"7fbd", x"7fbd", x"7fbe", x"7fbe", x"7fbe", 
    x"7fbe", x"7fbe", x"7fbf", x"7fbf", x"7fbf", x"7fbf", x"7fbf", x"7fc0", 
    x"7fc0", x"7fc0", x"7fc0", x"7fc0", x"7fc1", x"7fc1", x"7fc1", x"7fc1", 
    x"7fc1", x"7fc2", x"7fc2", x"7fc2", x"7fc2", x"7fc2", x"7fc2", x"7fc3", 
    x"7fc3", x"7fc3", x"7fc3", x"7fc3", x"7fc4", x"7fc4", x"7fc4", x"7fc4", 
    x"7fc4", x"7fc5", x"7fc5", x"7fc5", x"7fc5", x"7fc5", x"7fc6", x"7fc6", 
    x"7fc6", x"7fc6", x"7fc6", x"7fc6", x"7fc7", x"7fc7", x"7fc7", x"7fc7", 
    x"7fc7", x"7fc8", x"7fc8", x"7fc8", x"7fc8", x"7fc8", x"7fc8", x"7fc9", 
    x"7fc9", x"7fc9", x"7fc9", x"7fc9", x"7fca", x"7fca", x"7fca", x"7fca", 
    x"7fca", x"7fca", x"7fcb", x"7fcb", x"7fcb", x"7fcb", x"7fcb", x"7fcb", 
    x"7fcc", x"7fcc", x"7fcc", x"7fcc", x"7fcc", x"7fcd", x"7fcd", x"7fcd", 
    x"7fcd", x"7fcd", x"7fcd", x"7fce", x"7fce", x"7fce", x"7fce", x"7fce", 
    x"7fce", x"7fcf", x"7fcf", x"7fcf", x"7fcf", x"7fcf", x"7fcf", x"7fd0", 
    x"7fd0", x"7fd0", x"7fd0", x"7fd0", x"7fd0", x"7fd1", x"7fd1", x"7fd1", 
    x"7fd1", x"7fd1", x"7fd1", x"7fd2", x"7fd2", x"7fd2", x"7fd2", x"7fd2", 
    x"7fd2", x"7fd3", x"7fd3", x"7fd3", x"7fd3", x"7fd3", x"7fd3", x"7fd4", 
    x"7fd4", x"7fd4", x"7fd4", x"7fd4", x"7fd4", x"7fd5", x"7fd5", x"7fd5", 
    x"7fd5", x"7fd5", x"7fd5", x"7fd6", x"7fd6", x"7fd6", x"7fd6", x"7fd6", 
    x"7fd6", x"7fd6", x"7fd7", x"7fd7", x"7fd7", x"7fd7", x"7fd7", x"7fd7", 
    x"7fd8", x"7fd8", x"7fd8", x"7fd8", x"7fd8", x"7fd8", x"7fd8", x"7fd9", 
    x"7fd9", x"7fd9", x"7fd9", x"7fd9", x"7fd9", x"7fda", x"7fda", x"7fda", 
    x"7fda", x"7fda", x"7fda", x"7fda", x"7fdb", x"7fdb", x"7fdb", x"7fdb", 
    x"7fdb", x"7fdb", x"7fdb", x"7fdc", x"7fdc", x"7fdc", x"7fdc", x"7fdc", 
    x"7fdc", x"7fdc", x"7fdd", x"7fdd", x"7fdd", x"7fdd", x"7fdd", x"7fdd", 
    x"7fdd", x"7fde", x"7fde", x"7fde", x"7fde", x"7fde", x"7fde", x"7fde", 
    x"7fdf", x"7fdf", x"7fdf", x"7fdf", x"7fdf", x"7fdf", x"7fdf", x"7fe0", 
    x"7fe0", x"7fe0", x"7fe0", x"7fe0", x"7fe0", x"7fe0", x"7fe1", x"7fe1", 
    x"7fe1", x"7fe1", x"7fe1", x"7fe1", x"7fe1", x"7fe1", x"7fe2", x"7fe2", 
    x"7fe2", x"7fe2", x"7fe2", x"7fe2", x"7fe2", x"7fe3", x"7fe3", x"7fe3", 
    x"7fe3", x"7fe3", x"7fe3", x"7fe3", x"7fe3", x"7fe4", x"7fe4", x"7fe4", 
    x"7fe4", x"7fe4", x"7fe4", x"7fe4", x"7fe4", x"7fe5", x"7fe5", x"7fe5", 
    x"7fe5", x"7fe5", x"7fe5", x"7fe5", x"7fe5", x"7fe6", x"7fe6", x"7fe6", 
    x"7fe6", x"7fe6", x"7fe6", x"7fe6", x"7fe6", x"7fe7", x"7fe7", x"7fe7", 
    x"7fe7", x"7fe7", x"7fe7", x"7fe7", x"7fe7", x"7fe8", x"7fe8", x"7fe8", 
    x"7fe8", x"7fe8", x"7fe8", x"7fe8", x"7fe8", x"7fe8", x"7fe9", x"7fe9", 
    x"7fe9", x"7fe9", x"7fe9", x"7fe9", x"7fe9", x"7fe9", x"7fe9", x"7fea", 
    x"7fea", x"7fea", x"7fea", x"7fea", x"7fea", x"7fea", x"7fea", x"7fea", 
    x"7feb", x"7feb", x"7feb", x"7feb", x"7feb", x"7feb", x"7feb", x"7feb", 
    x"7feb", x"7fec", x"7fec", x"7fec", x"7fec", x"7fec", x"7fec", x"7fec", 
    x"7fec", x"7fec", x"7fed", x"7fed", x"7fed", x"7fed", x"7fed", x"7fed", 
    x"7fed", x"7fed", x"7fed", x"7fed", x"7fee", x"7fee", x"7fee", x"7fee", 
    x"7fee", x"7fee", x"7fee", x"7fee", x"7fee", x"7fef", x"7fef", x"7fef", 
    x"7fef", x"7fef", x"7fef", x"7fef", x"7fef", x"7fef", x"7fef", x"7fef", 
    x"7ff0", x"7ff0", x"7ff0", x"7ff0", x"7ff0", x"7ff0", x"7ff0", x"7ff0", 
    x"7ff0", x"7ff0", x"7ff1", x"7ff1", x"7ff1", x"7ff1", x"7ff1", x"7ff1", 
    x"7ff1", x"7ff1", x"7ff1", x"7ff1", x"7ff1", x"7ff2", x"7ff2", x"7ff2", 
    x"7ff2", x"7ff2", x"7ff2", x"7ff2", x"7ff2", x"7ff2", x"7ff2", x"7ff2", 
    x"7ff3", x"7ff3", x"7ff3", x"7ff3", x"7ff3", x"7ff3", x"7ff3", x"7ff3", 
    x"7ff3", x"7ff3", x"7ff3", x"7ff3", x"7ff4", x"7ff4", x"7ff4", x"7ff4", 
    x"7ff4", x"7ff4", x"7ff4", x"7ff4", x"7ff4", x"7ff4", x"7ff4", x"7ff4", 
    x"7ff5", x"7ff5", x"7ff5", x"7ff5", x"7ff5", x"7ff5", x"7ff5", x"7ff5", 
    x"7ff5", x"7ff5", x"7ff5", x"7ff5", x"7ff5", x"7ff6", x"7ff6", x"7ff6", 
    x"7ff6", x"7ff6", x"7ff6", x"7ff6", x"7ff6", x"7ff6", x"7ff6", x"7ff6", 
    x"7ff6", x"7ff6", x"7ff6", x"7ff7", x"7ff7", x"7ff7", x"7ff7", x"7ff7", 
    x"7ff7", x"7ff7", x"7ff7", x"7ff7", x"7ff7", x"7ff7", x"7ff7", x"7ff7", 
    x"7ff7", x"7ff8", x"7ff8", x"7ff8", x"7ff8", x"7ff8", x"7ff8", x"7ff8", 
    x"7ff8", x"7ff8", x"7ff8", x"7ff8", x"7ff8", x"7ff8", x"7ff8", x"7ff8", 
    x"7ff8", x"7ff9", x"7ff9", x"7ff9", x"7ff9", x"7ff9", x"7ff9", x"7ff9", 
    x"7ff9", x"7ff9", x"7ff9", x"7ff9", x"7ff9", x"7ff9", x"7ff9", x"7ff9", 
    x"7ff9", x"7ffa", x"7ffa", x"7ffa", x"7ffa", x"7ffa", x"7ffa", x"7ffa", 
    x"7ffa", x"7ffa", x"7ffa", x"7ffa", x"7ffa", x"7ffa", x"7ffa", x"7ffa", 
    x"7ffa", x"7ffa", x"7ffa", x"7ffa", x"7ffb", x"7ffb", x"7ffb", x"7ffb", 
    x"7ffb", x"7ffb", x"7ffb", x"7ffb", x"7ffb", x"7ffb", x"7ffb", x"7ffb", 
    x"7ffb", x"7ffb", x"7ffb", x"7ffb", x"7ffb", x"7ffb", x"7ffb", x"7ffb", 
    x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", 
    x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", 
    x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", 
    x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", 
    x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", 
    x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", 
    x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffe", x"7ffe", x"7ffe", 
    x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", 
    x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", 
    x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", 
    x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", 
    x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7fff", 
    x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", 
    x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", 
    x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", 
    x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", 
    x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", 
    x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", 
    x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff");

begin

PROCESS (CLK)
BEGIN
	if (rising_edge (clk)) then
		dsADD <= pdsADD;
		dcADD <= pdcADD;
		if ((sADD = x"4000") or (sADD = x"c000")) then
			sAz <= '1';
		else
			sAz <= '0';
		end if;
		if ((cADD = x"0000") or (cADD = x"8000")) then
			cAz <= '1';
		else
			cAz <= '0';
		end if;
		if (ADD(15 downto 14) = "00") then
			pdsADD <= '0';
			pdcADD <= '0';
			sADD <= "00" & ADD(13 downto 0);
			cADD <= "00" & (x"0" - ADD(13 downto 0));
		elsif (ADD(15 downto 14) = "01") then
			pdsADD <= '0';
			pdcADD <= '1';
			sADD <= "01" & (x"0" - ADD(13 downto 0));
			cADD <= "01" & ADD(13 downto 0);
		elsif (ADD(15 downto 14) = "10") then
			pdsADD <= '1';
			pdcADD <= '1';
			sADD <= "10" & ADD(13 downto 0);
			cADD <= "10" & (x"0" - ADD(13 downto 0));
		else -- (ADD(15 downto 14) = "11") then
			pdsADD <= '1';
			pdcADD <= '0';
			sADD <= "11" & (x"0" - ADD(13 downto 0));
			cADD <= "11" & ADD(13 downto 0);
		end if;
		msin <= isin(conv_integer(sADD(13 downto 0)));
		mcos <= isin(conv_integer(cADD(13 downto 0)));
		if (dsADD = '0') then
			if (sAz = '0') then
				nsin <= x"0" - msin;
			else
				nsin <= x"8001";
			end if;
		else
			if (sAz = '0') then
				nsin <= msin;
			else
				nsin <= x"7fff";
			end if;
			
		end if;
		if (dcADD = '0') then
			if (cAz = '0') then
				cos <= mcos;
			else
				cos <= x"7fff";
			end if;			
		else 
			if (cAz = '0') then
				cos <= x"0" - mcos;
			else
				cos <= x"8001";
			end if;
			
		end if;	
	end if;
END PROCESS;


end architecture;
