library IEEE;
use IEEE.std_logic_1164.all; 
use IEEE.std_logic_unsigned.all; 
use ieee.numeric_std.all;

entity bootloader_dp_32 is
  port (
    CLK:              in std_logic;
    WEA:  in std_logic;
    ENA:  in std_logic;
    MASKA:    in std_logic_vector(3 downto 0);
    ADDRA:         in std_logic_vector(11 downto 2);
    DIA:        in std_logic_vector(31 downto 0);
    DOA:         out std_logic_vector(31 downto 0);
    WEB:  in std_logic;
    ENB:  in std_logic;
    ADDRB:         in std_logic_vector(11 downto 2);
    DIB:        in std_logic_vector(31 downto 0);
    MASKB:    in std_logic_vector(3 downto 0);
    DOB:         out std_logic_vector(31 downto 0)
  );
end entity bootloader_dp_32;

architecture behave of bootloader_dp_32 is

  subtype RAM_WORD is STD_LOGIC_VECTOR (31 downto 0);
  type RAM_TABLE is array (0 to 1023) of RAM_WORD;
 shared variable RAM: RAM_TABLE := RAM_TABLE'(
x"0b0b0b94",x"d5040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b94",x"f1040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fd0608",x"72830609",x"81058205",x"832b2a83",x"ffff0652",x"04000000",x"00000000",x"00000000",x"71fd0608",x"83ffff73",x"83060981",x"05820583",x"2b2b0906",x"7383ffff",x"0b0b0b0b",x"83a70400",x"72098105",x"72057373",x"09060906",x"73097306",x"070a8106",x"53510400",x"00000000",x"00000000",x"72722473",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71737109",x"71068106",x"30720a10",x"0a720a10",x"0a31050a",x"81065151",x"53510400",x"00000000",x"72722673",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"c3040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"720a722b",x"0a535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72729f06",x"0981050b",x"0b0b88a6",x"05040000",x"00000000",x"00000000",x"00000000",x"00000000",x"72722aff",x"739f062a",x"0974090a",x"8106ff05",x"06075351",x"04000000",x"00000000",x"00000000",x"71715351",x"020d0406",x"73830609",x"81058205",x"832b0b2b",x"0772fc06",x"0c515104",x"00000000",x"72098105",x"72050970",x"81050906",x"0a810653",x"51040000",x"00000000",x"00000000",x"00000000",x"72098105",x"72050970",x"81050906",x"0a098106",x"53510400",x"00000000",x"00000000",x"00000000",x"71098105",x"52040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72720981",x"05055351",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097206",x"73730906",x"07535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fc0608",x"72830609",x"81058305",x"1010102a",x"81ff0652",x"04000000",x"00000000",x"00000000",x"71fc0608",x"0b0b0b97",x"88738306",x"10100508",x"060b0b0b",x"88a90400",x"00000000",x"00000000",x"0b0b0b88",x"f7040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"df040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097081",x"0509060a",x"8106ff05",x"70547106",x"73097274",x"05ff0506",x"07515151",x"04000000",x"72097081",x"0509060a",x"098106ff",x"05705471",x"06730972",x"7405ff05",x"06075151",x"51040000",x"05ff0504",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"810b0b0b",x"0b9aac0c",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71810552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"02840572",x"10100552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"717105ff",x"05715351",x"020d0400",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"81d43f8e",x"d73f0410",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10105351",x"047381ff",x"06738306",x"09810583",x"05101010",x"2b0772fc",x"060c5151",x"043c0472",x"72807281",x"06ff0509",x"72060571",x"1052720a",x"100a5372",x"ed385151",x"53510488",x"088c0890",x"08757595",x"c72d5050",x"88085690",x"0c8c0c88",x"0c510488",x"088c0890",x"08757595",x"832d5050",x"88085690",x"0c8c0c88",x"0c510488",x"088c0890",x"088dee2d",x"900c8c0c",x"880c04ff",x"3d0d0b0b",x"0b9abc33",x"5170a638",x"9ab80870",x"08525270",x"802e9238",x"84129ab8",x"0c702d9a",x"b8087008",x"525270f0",x"38810b0b",x"0b0b9abc",x"34833d0d",x"0404803d",x"0d0b0b0b",x"9ae00880",x"2e8e380b",x"0b0b0b80",x"0b802e09",x"81068538",x"823d0d04",x"0b0b0b9a",x"e0510b0b",x"0bf6813f",x"823d0d04",x"04ff3d0d",x"80c48080",x"84527108",x"70822a70",x"81065151",x"5170f338",x"833d0d04",x"ff3d0d80",x"c4808084",x"52710870",x"812a7081",x"06515151",x"70f33873",x"82900a0c",x"833d0d04",x"ff3d0d73",x"8f065289",x"72278738",x"80d71251",x"8439b012",x"518aa02d",x"833d0d04",x"fd3d0d75",x"54733370",x"81ff0653",x"5371802e",x"8e387281",x"ff06518a",x"a02d8114",x"54e73985",x"3d0d04ff",x"3d0d7370",x"842a5252",x"8ac02d71",x"518ac02d",x"833d0d04",x"ff3d0d73",x"70982a52",x"528aff2d",x"71902a51",x"8aff2d71",x"882a518a",x"ff2d7151",x"8aff2d83",x"3d0d04ff",x"3d0d7370",x"08515180",x"c8808084",x"70087084",x"80800772",x"0c525283",x"3d0d04ff",x"3d0d80c8",x"80808470",x"0870fbff",x"ff06720c",x"5252833d",x"0d04a090",x"0ba0800c",x"9ac00ba0",x"840c94ea",x"2dff3d0d",x"73518b71",x"0c901152",x"98808072",x"0c80720c",x"700883ff",x"ff06880c",x"833d0d04",x"fa3d0d78",x"7a7dff1e",x"57575853",x"73ff2ea7",x"38805684",x"5275730c",x"72088818",x"0cff1252",x"71f33874",x"84167408",x"720cff16",x"56565273",x"ff2e0981",x"06dd3888",x"3d0d04f8",x"3d0d80c0",x"80808457",x"83d00a59",x"8bd32d76",x"518bf92d",x"9ac07088",x"08101098",x"80840571",x"70840553",x"0c5656fb",x"8084a1ad",x"750c9798",x"0b88170c",x"8070780c",x"770c7608",x"83ffff06",x"569fdf80",x"0b880827",x"8338ff39",x"83ffff79",x"0ca08054",x"88085378",x"5276518c",x"982d7651",x"8bb72d78",x"08557476",x"2e893880",x"c3518aa0",x"2dff39a0",x"84085574",x"faa094a6",x"802e8938",x"80c2518a",x"a02dff39",x"900a7008",x"70ffbf06",x"720c5656",x"8a852d8b",x"ea2dff3d",x"0d9acc08",x"81119acc",x"0c518390",x"0a700870",x"feff0672",x"0c525283",x"3d0d04ff",x"b23d0d84",x"80b30b80",x"c4808084",x"0c80c880",x"80a453fb",x"ffff7308",x"70720675",x"0c535480",x"c8808094",x"70087076",x"06720c53",x"53800b80",x"fc8097a8",x"52568adc",x"2d80fc80",x"97cc518a",x"dc2d7553",x"fad5aad5",x"aa70740c",x"73085354",x"71742e09",x"810681f8",x"3885aad5",x"aad57074",x"0c730853",x"5471742e",x"09810681",x"e338faaa",x"eacada70",x"740c7308",x"53547174",x"2e098106",x"81ce3885",x"d7c1d68f",x"70740c73",x"08535471",x"742e0981",x"0681b938",x"8070740c",x"73085354",x"71742e09",x"810681a8",x"38ff7074",x"0c730853",x"5471742e",x"09810681",x"973880d5",x"0a70740c",x"73085354",x"71742e09",x"81068184",x"3885a880",x"8070740c",x"73085354",x"71742e09",x"810680f0",x"3882d480",x"70740c73",x"08535471",x"742e0981",x"0680dd38",x"81aa7074",x"0c730853",x"5471742e",x"09810680",x"cb388413",x"53728880",x"802e0981",x"06feb138",x"75802e80",x"c03880fc",x"8097ec51",x"8adc2d72",x"518b942d",x"80fc8098",x"80518adc",x"2d73518b",x"942d80fc",x"80988c51",x"8adc2d71",x"518b942d",x"80fc8097",x"c8518adc",x"2d83f839",x"8156c139",x"815680ca",x"3980fc80",x"989c518a",x"dc2d80fc",x"8098b451",x"8adc2d75",x"76545473",x"73708405",x"550c8114",x"54728880",x"802e0981",x"06ed3880",x"70555372",x"08527174",x"2e098106",x"c3388114",x"84145454",x"72888080",x"2e098106",x"e6387580",x"2ea03880",x"fc8097ec",x"518adc2d",x"72518b94",x"2d80fc80",x"97c8518a",x"dc2d8387",x"39815680",x"d53980fc",x"8098d451",x"8adc2d80",x"fc8098f4",x"518adc2d",x"75765654",x"73757081",x"05573481",x"145474a0",x"80802e09",x"8106ed38",x"80705555",x"74337081",x"ff067581",x"ff065551",x"5271732e",x"098106ff",x"b8388114",x"81165654",x"74a08080",x"2e098106",x"db387580",x"2ea03880",x"fc80999c",x"518adc2d",x"74518b94",x"2d80fc80",x"97c8518a",x"dc2d828f",x"39815681",x"c73980fc",x"8099b451",x"8adc2d80",x"fc8099d4",x"518adc2d",x"7553fad5",x"aad5aa54",x"7274740c",x"73085355",x"71742e09",x"8106d238",x"80d57334",x"85adaad5",x"aa730853",x"5771772e",x"098106ff",x"bc388113",x"74740c73",x"08535571",x"742e0981",x"06ffaa38",x"80d57534",x"fad2d6d5",x"aa730853",x"5771772e",x"098106ff",x"94388115",x"74740c73",x"08535571",x"742e0981",x"06ff8238",x"80d57534",x"fad5a9ab",x"aa730853",x"5771772e",x"098106fe",x"ec388115",x"74740c73",x"08535571",x"742e0981",x"06feda38",x"80d57534",x"fad5aad4",x"d5730853",x"5771772e",x"098106fe",x"c4388413",x"53728880",x"802e0981",x"06fed538",x"75802eb6",x"3880fc80",x"999c518a",x"dc2d7451",x"8b942d80",x"fc8099f8",x"518adc2d",x"76518b94",x"2d80fc80",x"988c518a",x"dc2d7151",x"8b942d80",x"fc8097c8",x"518adc2d",x"8a3980fc",x"809a8851",x"8adc2dff",x"39ff3d0d",x"80528051",x"8e8b2d83",x"3d0d049f",x"fff80d8c",x"d3049fff",x"f80da088",x"0488088c",x"08a0802d",x"8c0c880c",x"810b80d0",x"0a0c04fb",x"3d0d7779",x"55558056",x"757524ab",x"38807424",x"9d388053",x"73527451",x"80e13f88",x"08547580",x"2e853888",x"08305473",x"880c873d",x"0d047330",x"76813257",x"54dc3974",x"30558156",x"738025d2",x"38ec39fa",x"3d0d787a",x"57558057",x"767524a4",x"38759f2c",x"54815375",x"74327431",x"5274519b",x"3f880854",x"76802e85",x"38880830",x"5473880c",x"883d0d04",x"74305581",x"57d739fc",x"3d0d7678",x"53548153",x"80747326",x"52557280",x"2e983870",x"802ea938",x"807224a4",x"38711073",x"10757226",x"53545272",x"ea387351",x"78833874",x"5170880c",x"863d0d04",x"72812a72",x"812a5353",x"72802ee6",x"38717426",x"ef387372",x"31757407",x"74812a74",x"812a5555",x"5654e539",x"ff3d0d9a",x"d40bfc05",x"70085252",x"70ff2e91",x"38702dfc",x"12700852",x"5270ff2e",x"098106f1",x"38833d0d",x"0404f29b",x"3f040000",x"00ffffff",x"ff00ffff",x"ffff00ff",x"ffffff00",x"01090600",x"0007ef80",x"05b8d800",x"a4051300",x"5a505569",x"6e6f204d",x"656d6f72",x"79205465",x"73746572",x"20737461",x"7274696e",x"672e0d0a",x"0d0a0000",x"53746172",x"74696e67",x"2073696d",x"706c6520",x"70617474",x"65726e20",x"74657374",x"2e2e2e00",x"4572726f",x"72206174",x"20616464",x"72657373",x"20307800",x"3a207772",x"6f746520",x"30780000",x"2c207265",x"61642062",x"61636b20",x"30780000",x"53746570",x"20312028",x"776f7264",x"29207061",x"73736564",x"2e0d0a00",x"53746172",x"74696e67",x"20696e63",x"72656d65",x"6e74616c",x"20746573",x"742e2e2e",x"00000000",x"53746570",x"20322028",x"696e6372",x"656d656e",x"74616c29",x"20706173",x"7365642e",x"0d0a0000",x"53746172",x"74696e67",x"20627974",x"65776973",x"6520696e",x"6372656d",x"656e7461",x"6c207465",x"73742e2e",x"2e000000",x"0d0a4572",x"726f7220",x"61742061",x"64647265",x"73732030",x"78000000",x"53746570",x"20332028",x"62797465",x"2d776973",x"65292070",x"61737365",x"642e0d0a",x"00000000",x"53746172",x"74696e67",x"20656e64",x"69616e20",x"62797465",x"2d776973",x"65207465",x"73742e2e",x"2e000000",x"3a206578",x"70656374",x"65642030",x"78000000",x"53746570",x"20342028",x"656e6469",x"616e2062",x"7974652d",x"77697365",x"29207061",x"73736564",x"2e0d0a00",x"00000000",x"00000000",x"00000000",x"00000d5c",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"ffffffff",x"00000000",x"ffffffff",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000");

begin

  process (clk)
  begin
    if rising_edge(clk) then
      if ENA='1' then
        if WEA='1' then
          RAM(conv_integer(ADDRA) ) := DIA;
        end if;
        DOA <= RAM(conv_integer(ADDRA)) ;
      end if;
    end if;
  end process;  

  process (clk)
  begin
    if rising_edge(clk) then
      if ENB='1' then
        if WEB='1' then
          RAM( conv_integer(ADDRB) ) := DIB;
        end if;
        DOB <= RAM(conv_integer(ADDRB)) ;
      end if;
    end if;
  end process;  
end behave;
