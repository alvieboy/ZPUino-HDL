library IEEE;
use IEEE.std_logic_1164.all; 
use IEEE.std_logic_unsigned.all; 
use ieee.numeric_std.all;

entity bootloader_dp_32 is
  port (
    CLK:              in std_logic;
    WEA:  in std_logic;
    ENA:  in std_logic;
    MASKA:    in std_logic_vector(3 downto 0);
    ADDRA:         in std_logic_vector(11 downto 2);
    DIA:        in std_logic_vector(31 downto 0);
    DOA:         out std_logic_vector(31 downto 0);
    WEB:  in std_logic;
    ENB:  in std_logic;
    ADDRB:         in std_logic_vector(11 downto 2);
    DIB:        in std_logic_vector(31 downto 0);
    MASKB:    in std_logic_vector(3 downto 0);
    DOB:         out std_logic_vector(31 downto 0)
  );
end entity bootloader_dp_32;

architecture behave of bootloader_dp_32 is

  subtype RAM_WORD is STD_LOGIC_VECTOR (31 downto 0);
  type RAM_TABLE is array (0 to 1023) of RAM_WORD;
 shared variable RAM: RAM_TABLE := RAM_TABLE'(
x"0b0b0b97",x"82040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b96",x"ed040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fd0608",x"72830609",x"81058205",x"832b2a83",x"ffff0652",x"04000000",x"00000000",x"00000000",x"71fd0608",x"83ffff73",x"83060981",x"05820583",x"2b2b0906",x"7383ffff",x"0b0b0b0b",x"83a70400",x"72098105",x"72057373",x"09060906",x"73097306",x"070a8106",x"53510400",x"00000000",x"00000000",x"72722473",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71737109",x"71068106",x"30720a10",x"0a720a10",x"0a31050a",x"81065151",x"53510400",x"00000000",x"72722673",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"cc040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"720a722b",x"0a535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72729f06",x"0981050b",x"0b0b88af",x"05040000",x"00000000",x"00000000",x"00000000",x"00000000",x"72722aff",x"739f062a",x"0974090a",x"8106ff05",x"06075351",x"04000000",x"00000000",x"00000000",x"71715351",x"020d0406",x"73830609",x"81058205",x"832b0b2b",x"0772fc06",x"0c515104",x"00000000",x"72098105",x"72050970",x"81050906",x"0a810653",x"51040000",x"00000000",x"00000000",x"00000000",x"72098105",x"72050970",x"81050906",x"0a098106",x"53510400",x"00000000",x"00000000",x"00000000",x"71098105",x"52040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72720981",x"05055351",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097206",x"73730906",x"07535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fc0608",x"72830609",x"81058305",x"1010102a",x"81ff0652",x"04000000",x"00000000",x"00000000",x"71fc0608",x"0b0b0b99",x"ec738306",x"10100508",x"060b0b0b",x"88b20400",x"00000000",x"00000000",x"0b0b0b89",x"80040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"e8040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097081",x"0509060a",x"8106ff05",x"70547106",x"73097274",x"05ff0506",x"07515151",x"04000000",x"72097081",x"0509060a",x"098106ff",x"05705471",x"06730972",x"7405ff05",x"06075151",x"51040000",x"05ff0504",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"810b0b0b",x"0b9aa40c",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71810552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"02840572",x"10100552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"717105ff",x"05715351",x"020d0400",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"81dd3f91",x"bd3f0400",x"00000000",x"00000000",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101053",x"51047381",x"ff067383",x"06098105",x"83051010",x"102b0772",x"fc060c51",x"51043c04",x"72728072",x"8106ff05",x"09720605",x"71105272",x"0a100a53",x"72ed3851",x"51535104",x"88088c08",x"90087575",x"98ad2d50",x"50880856",x"900c8c0c",x"880c5104",x"88088c08",x"90087575",x"97e92d50",x"50880856",x"900c8c0c",x"880c5104",x"88088c08",x"90088df6",x"2d900c8c",x"0c880c04",x"ff3d0d0b",x"0b0b9ac8",x"335170a6",x"389ab008",x"70085252",x"70802e92",x"3884129a",x"b00c702d",x"9ab00870",x"08525270",x"f038810b",x"0b0b0b9a",x"c834833d",x"0d040480",x"3d0d0b0b",x"0b9af408",x"802e8e38",x"0b0b0b0b",x"800b802e",x"09810685",x"38823d0d",x"040b0b0b",x"9af4510b",x"0b0bf5f8",x"3f823d0d",x"0404ff3d",x"0d80c480",x"80845271",x"0870822a",x"70810651",x"515170f3",x"38833d0d",x"04ff3d0d",x"80c48080",x"84527108",x"70812a70",x"81065151",x"5170f338",x"7382900a",x"0c833d0d",x"04fe3d0d",x"747080dc",x"8080880c",x"7081ff06",x"ff831154",x"51537181",x"268d3880",x"fd518aa9",x"2d72a032",x"51833972",x"518aa92d",x"843d0d04",x"803d0d83",x"ffff0b83",x"d00a0c80",x"fe518aa9",x"2d823d0d",x"04ff3d0d",x"83d00a08",x"70882a52",x"528ac92d",x"7181ff06",x"518ac92d",x"80fe518a",x"a92d833d",x"0d048386",x"cf0b80cc",x"8080880c",x"800b80cc",x"8080840c",x"9f0b8390",x"0a0c04ff",x"3d0d7370",x"08515180",x"c8808084",x"70087084",x"80800772",x"0c525283",x"3d0d04ff",x"3d0d80c8",x"80808470",x"0870fbff",x"ff06720c",x"5252833d",x"0d04a090",x"0ba0800c",x"9acc0ba0",x"840c96e5",x"2dff3d0d",x"73518b71",x"0c901152",x"98808072",x"0c80720c",x"700883ff",x"ff06880c",x"833d0d04",x"fa3d0d78",x"7a7dff1e",x"57575853",x"73ff2ea7",x"38805684",x"5275730c",x"72088818",x"0cff1252",x"71f33874",x"84167408",x"720cff16",x"56565273",x"ff2e0981",x"06dd3888",x"3d0d04f9",x"3d0d80d0",x"80808456",x"83d00a58",x"8be32d75",x"518c892d",x"9acc7088",x"08101098",x"80840571",x"70840553",x"0c5657fb",x"8084a1ad",x"750c9ab4",x"0b88180c",x"8070770c",x"760c7508",x"7083ffff",x"06515783",x"ffff780c",x"a0805488",x"08537752",x"75518ca8",x"2d75518b",x"c72d7708",x"5574772e",x"893880c3",x"518aa92d",x"ff39a084",x"085574fb",x"d888b480",x"2e893880",x"c2518aa9",x"2dff3980",x"d00a7008",x"70ffbf06",x"720c5656",x"8a8e2d8b",x"fa2dff3d",x"0d9ad808",x"81119ad8",x"0c518390",x"0a700870",x"feff0672",x"0c525283",x"3d0d0480",x"3d0d8af8",x"2d728180",x"07518ac9",x"2d8b8d2d",x"823d0d04",x"fe3d0d80",x"d0808084",x"538be32d",x"85730c80",x"730c7208",x"7081ff06",x"74535152",x"8bc72d71",x"880c843d",x"0d04fc3d",x"0d768111",x"33821233",x"7181800a",x"29718480",x"80290583",x"14337082",x"80291284",x"16335271",x"05a08005",x"86168517",x"33575253",x"53555755",x"53ff1353",x"72ff2e91",x"38737081",x"05553352",x"71757081",x"055734e9",x"3989518e",x"932d863d",x"0d04f93d",x"0d795780",x"d0808084",x"568be32d",x"81173382",x"18337182",x"80290553",x"5371802e",x"94388517",x"72555372",x"70810554",x"33760cff",x"145473f3",x"38831733",x"84183371",x"82802905",x"56528054",x"73752797",x"38735877",x"760c7317",x"76085353",x"71733481",x"14547474",x"26ed3875",x"518bc72d",x"8af82d81",x"84518ac9",x"2d74882a",x"518ac92d",x"74518ac9",x"2d805473",x"75278f38",x"73177033",x"52528ac9",x"2d811454",x"ee398b8d",x"2d893d0d",x"0404fc3d",x"0d768111",x"33821233",x"71902b71",x"882b0783",x"14337072",x"07882b84",x"16337107",x"51525357",x"57545288",x"518e932d",x"81ff518a",x"a92d80c4",x"80808453",x"72087081",x"2a708106",x"51515271",x"f3387384",x"80800780",x"c4808084",x"0c863d0d",x"04fe3d0d",x"8ea82d88",x"08880881",x"06535371",x"f3388af8",x"2d818351",x"8ac92d72",x"518ac92d",x"8b8d2d84",x"3d0d04fe",x"3d0d800b",x"9ad80c8a",x"f82d8181",x"518ac92d",x"9ab45393",x"52727081",x"05543351",x"8ac92dff",x"125271ff",x"2e098106",x"ec388b8d",x"2d843d0d",x"04fe3d0d",x"800b9ad8",x"0c8af82d",x"8182518a",x"c92d80d0",x"80808452",x"8be32d81",x"f90a0b80",x"d080809c",x"0c710872",x"52538bc7",x"2d729ae0",x"0c72902a",x"518ac92d",x"9ae00888",x"2a518ac9",x"2d9ae008",x"518ac92d",x"8ea82d88",x"08518ac9",x"2d8b8d2d",x"843d0d04",x"803d0d81",x"0b9adc0c",x"800b8390",x"0a0c8551",x"8e932d82",x"3d0d0480",x"3d0d800b",x"9adc0c8b",x"ae2d8651",x"8e932d82",x"3d0d04fd",x"3d0d80d0",x"80808454",x"8a518e93",x"2d8be32d",x"9acc7452",x"538c892d",x"72880810",x"10988084",x"05717084",x"05530c52",x"fb8084a1",x"ad720c9a",x"b40b8814",x"0c73518b",x"c72d8a8e",x"2d8bfa2d",x"ffab3d0d",x"80d93d08",x"56800b9a",x"dc0c800b",x"9ad80c80",x"0bdf8017",x"9ab97190",x"2a715656",x"57555772",x"72708105",x"54347388",x"2a537272",x"34738216",x"34758b16",x"348df60b",x"a0800c80",x"c4808084",x"558480b5",x"750c80c8",x"8080a453",x"fbffff73",x"08707206",x"750c5354",x"80c88080",x"94700870",x"7606720c",x"5353880b",x"80c08080",x"840c900a",x"5381730c",x"8bae2dfe",x"88880b80",x"dc808084",x"0c81f20b",x"80d00a0c",x"80d08080",x"84705252",x"8bc72d8b",x"e32d7151",x"8bc72d76",x"77767593",x"3d41415b",x"5b5b83d0",x"0a5c7808",x"70810651",x"52719d38",x"9adc0853",x"72f0389a",x"d8085287",x"e87227e6",x"38727e0c",x"7283900a",x"0c96dd2d",x"82900a08",x"5379802e",x"81b43872",x"80fe2e09",x"810680f4",x"3876802e",x"c138807d",x"7857575a",x"827727ff",x"b53883ff",x"ff7c0c79",x"fe185353",x"79722798",x"3880dc80",x"80887255",x"58721670",x"33790c52",x"81135373",x"7326f238",x"ff157611",x"547605ff",x"05703374",x"33707288",x"2b077f08",x"53515551",x"5271732e",x"098106fe",x"ed387533",x"53728a26",x"fee43872",x"101099f8",x"05765270",x"08515271",x"2dfed339",x"7280fd2e",x"09810686",x"38815bfe",x"c5397682",x"9f269e38",x"7a802e87",x"388073a0",x"32545b80",x"d73d7705",x"fde00552",x"72723481",x"1757fea2",x"39805afe",x"9d397280",x"fe2e0981",x"06fe9338",x"7957ff7c",x"0c81775c",x"5afe8739",x"ff3d0d97",x"bd2d7352",x"805193a4",x"2d833d0d",x"049fffff",x"f80d8ce3",x"049fffff",x"f80da088",x"04880880",x"c0808088",x"08a08008",x"2d50880c",x"810b900a",x"0c048070",x"0cfaad95",x"b4da0b81",x"80807171",x"0c718008",x"2e873870",x"1151978e",x"045196cc",x"2d000000",x"00000000",x"00000000",x"00000000",x"820b80c0",x"8080900c",x"0b0b0b04",x"0083f00a",x"0b800ba0",x"80721208",x"720c8412",x"5271712e",x"ff05f238",x"028c050d",x"97b00400",x"00000000",x"00000000",x"00000000",x"00fb3d0d",x"77795555",x"80567575",x"24ab3880",x"74249d38",x"80537352",x"745180e1",x"3f880854",x"75802e85",x"38880830",x"5473880c",x"873d0d04",x"73307681",x"325754dc",x"39743055",x"81567380",x"25d238ec",x"39fa3d0d",x"787a5755",x"80577675",x"24a43875",x"9f2c5481",x"53757432",x"74315274",x"519b3f88",x"08547680",x"2e853888",x"08305473",x"880c883d",x"0d047430",x"558157d7",x"39fc3d0d",x"76785354",x"81538074",x"73265255",x"72802e98",x"3870802e",x"a9388072",x"24a43871",x"10731075",x"72265354",x"5272ea38",x"73517883",x"38745170",x"880c863d",x"0d047281",x"2a72812a",x"53537280",x"2ee63871",x"7426ef38",x"73723175",x"74077481",x"2a74812a",x"55555654",x"e539ff3d",x"0d9ae80b",x"fc057008",x"525270ff",x"2e913870",x"2dfc1270",x"08525270",x"ff2e0981",x"06f13883",x"3d0d0404",x"efbe3f04",x"00ffffff",x"ff00ffff",x"ffff00ff",x"ffffff00",x"000008af",x"000008e1",x"00000889",x"000007a2",x"00000938",x"0000094f",x"00000835",x"00000836",x"0000074e",x"00000963",x"00000000",x"00000000",x"00000000",x"00000d70",x"01090600",x"00000000",x"05f5e100",x"bb021a00",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"ffffffff",x"00000000",x"ffffffff",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000");

begin

  process (clk)
  begin
    if rising_edge(clk) then
      if ENA='1' then
        if WEA='1' then
          RAM(conv_integer(ADDRA) ) := DIA;
        end if;
        DOA <= RAM(conv_integer(ADDRA)) ;
      end if;
    end if;
  end process;  

  process (clk)
  begin
    if rising_edge(clk) then
      if ENB='1' then
        if WEB='1' then
          RAM( conv_integer(ADDRB) ) := DIB;
        end if;
        DOB <= RAM(conv_integer(ADDRB)) ;
      end if;
    end if;
  end process;  
end behave;
