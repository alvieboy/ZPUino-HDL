library IEEE;
use IEEE.std_logic_1164.all; 
use IEEE.std_logic_unsigned.all; 
use ieee.numeric_std.all;

entity bootloader_dp_32 is
  port (
    CLK:              in std_logic;
    WEA:  in std_logic;
    ENA:  in std_logic;
    MASKA:    in std_logic_vector(3 downto 0);
    ADDRA:         in std_logic_vector(11 downto 2);
    DIA:        in std_logic_vector(31 downto 0);
    DOA:         out std_logic_vector(31 downto 0);
    WEB:  in std_logic;
    ENB:  in std_logic;
    ADDRB:         in std_logic_vector(11 downto 2);
    DIB:        in std_logic_vector(31 downto 0);
    MASKB:    in std_logic_vector(3 downto 0);
    DOB:         out std_logic_vector(31 downto 0)
  );
end entity bootloader_dp_32;

architecture behave of bootloader_dp_32 is

  subtype RAM_WORD is STD_LOGIC_VECTOR (31 downto 0);
  type RAM_TABLE is array (0 to 1023) of RAM_WORD;
 shared variable RAM: RAM_TABLE := RAM_TABLE'(
x"0b0b0b97",x"95040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b97",x"b6040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fd0608",x"72830609",x"81058205",x"832b2a83",x"ffff0652",x"04000000",x"00000000",x"00000000",x"71fd0608",x"83ffff73",x"83060981",x"05820583",x"2b2b0906",x"7383ffff",x"0b0b0b0b",x"83a70400",x"72098105",x"72057373",x"09060906",x"73097306",x"070a8106",x"53510400",x"00000000",x"00000000",x"72722473",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71737109",x"71068106",x"30720a10",x"0a720a10",x"0a31050a",x"81065151",x"53510400",x"00000000",x"72722673",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"cc040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"720a722b",x"0a535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72729f06",x"0981050b",x"0b0b88af",x"05040000",x"00000000",x"00000000",x"00000000",x"00000000",x"72722aff",x"739f062a",x"0974090a",x"8106ff05",x"06075351",x"04000000",x"00000000",x"00000000",x"71715351",x"020d0406",x"73830609",x"81058205",x"832b0b2b",x"0772fc06",x"0c515104",x"00000000",x"72098105",x"72050970",x"81050906",x"0a810653",x"51040000",x"00000000",x"00000000",x"00000000",x"72098105",x"72050970",x"81050906",x"0a098106",x"53510400",x"00000000",x"00000000",x"00000000",x"71098105",x"52040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72720981",x"05055351",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097206",x"73730906",x"07535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fc0608",x"72830609",x"81058305",x"1010102a",x"81ff0652",x"04000000",x"00000000",x"00000000",x"71fc0608",x"0b0b0b9d",x"cc738306",x"10100508",x"060b0b0b",x"88b20400",x"00000000",x"00000000",x"0b0b0b89",x"80040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"e8040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097081",x"0509060a",x"8106ff05",x"70547106",x"73097274",x"05ff0506",x"07515151",x"04000000",x"72097081",x"0509060a",x"098106ff",x"05705471",x"06730972",x"7405ff05",x"06075151",x"51040000",x"05ff0504",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"810b0b0b",x"0b9e940c",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71810552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"02840572",x"10100552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"717105ff",x"05715351",x"020d0400",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"81dd3f95",x"9a3f0400",x"00000000",x"00000000",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101053",x"51047381",x"ff067383",x"06098105",x"83051010",x"102b0772",x"fc060c51",x"51043c04",x"72728072",x"8106ff05",x"09720605",x"71105272",x"0a100a53",x"72ed3851",x"51535104",x"88088c08",x"90087575",x"98cd2d50",x"50880856",x"900c8c0c",x"880c5104",x"88088c08",x"90087575",x"98892d50",x"50880856",x"900c8c0c",x"880c5104",x"88088c08",x"90088e8d",x"2d900c8c",x"0c880c04",x"ff3d0d0b",x"0b0b9ea4",x"335170a6",x"389ea008",x"70085252",x"70802e92",x"3884129e",x"a00c702d",x"9ea00870",x"08525270",x"f038810b",x"0b0b0b9e",x"a434833d",x"0d040480",x"3d0d0b0b",x"0b9ed008",x"802e8e38",x"0b0b0b0b",x"800b802e",x"09810685",x"38823d0d",x"040b0b0b",x"9ed0510b",x"0b0bf5f8",x"3f823d0d",x"0404ff3d",x"0d80c480",x"80845271",x"0870822a",x"70810651",x"515170f3",x"38833d0d",x"04ff3d0d",x"80c48080",x"84527108",x"70812a70",x"81065151",x"5170f338",x"7382900a",x"0c833d0d",x"04fe3d0d",x"747080dc",x"8080880c",x"7081ff06",x"ff831154",x"51537181",x"268d3880",x"fd518aa9",x"2d72a032",x"51833972",x"518aa92d",x"843d0d04",x"803d0d83",x"ffff0b83",x"d00a0c80",x"fe518aa9",x"2d823d0d",x"04ff3d0d",x"83d00a08",x"70882a52",x"528ac92d",x"7181ff06",x"518ac92d",x"80fe518a",x"a92d833d",x"0d048386",x"cf0b80cc",x"8080880c",x"800b80cc",x"8080840c",x"9f0b8390",x"0a0c8e8d",x"0ba0800c",x"810b900a",x"0c04ff3d",x"0d737008",x"515180c8",x"80808470",x"08708480",x"8007720c",x"5252833d",x"0d04ff3d",x"0d80c880",x"80847008",x"70fbffff",x"06720c52",x"52833d0d",x"04a0900b",x"a0800c9e",x"a80ba084",x"0c97ae2d",x"ff3d0d73",x"518b710c",x"90115280",x"dc808072",x"0c80720c",x"700883ff",x"ff06880c",x"833d0d04",x"fa3d0d78",x"7a7dff1e",x"57575853",x"73ff2ea7",x"38805684",x"5275730c",x"72088818",x"0cff1252",x"71f33874",x"84167408",x"720cff16",x"56565273",x"ff2e0981",x"06dd3888",x"3d0d04f8",x"3d0d80d0",x"80808457",x"83d00a59",x"8bee2d76",x"518c942d",x"9ea87088",x"08101080",x"dc808405",x"71708405",x"530c5656",x"fb8084a1",x"ad750c9e",x"840b8817",x"0c807078",x"0c770c76",x"0883ffff",x"06569fff",x"df800b88",x"08278338",x"ff3983ff",x"ff790ca0",x"80548808",x"53785276",x"518cb42d",x"76518bd2",x"2d780855",x"74762e89",x"3880c351",x"8aa92dff",x"39a08408",x"5574fbd0",x"84b4802e",x"893880c2",x"518aa92d",x"ff3980d0",x"0a700870",x"ffbf0672",x"0c56568a",x"8e2d8c85",x"2dff3d0d",x"9eb40881",x"119eb40c",x"5183900a",x"700870fe",x"ff06720c",x"5252833d",x"0d04803d",x"0d8af82d",x"72818007",x"518ac92d",x"8b8d2d82",x"3d0d04fe",x"3d0d80d0",x"80808453",x"8bee2d85",x"730c8073",x"0c720870",x"81ff0674",x"5351528b",x"d22d7188",x"0c843d0d",x"04fc3d0d",x"76811133",x"82123371",x"81800a29",x"71848080",x"29058314",x"33708280",x"29128416",x"33527105",x"a0800586",x"16851733",x"57525353",x"55575553",x"ff135372",x"ff2e9138",x"73708105",x"55335271",x"75708105",x"5734e939",x"89518eaa",x"2d863d0d",x"04f93d0d",x"795780d0",x"80808456",x"8bee2d81",x"17338218",x"33718280",x"29055353",x"71802e94",x"38851772",x"55537270",x"81055433",x"760cff14",x"5473f338",x"83173384",x"18337182",x"80290556",x"52805473",x"75279738",x"73587776",x"0c731776",x"08535371",x"73348114",x"54747426",x"ed387551",x"8bd22d8a",x"f82d8184",x"518ac92d",x"74882a51",x"8ac92d74",x"518ac92d",x"80547375",x"278f3873",x"17703352",x"528ac92d",x"811454ee",x"398b8d2d",x"893d0d04",x"04fc3d0d",x"76811133",x"82123371",x"902b7188",x"2b078314",x"33707207",x"882b8416",x"33710751",x"52535757",x"54528851",x"8eaa2d81",x"ff518aa9",x"2d80c480",x"80845372",x"0870812a",x"70810651",x"515271f3",x"38738480",x"800780c4",x"8080840c",x"863d0d04",x"fe3d0d8e",x"bf2d8808",x"88088106",x"535371f3",x"388af82d",x"8183518a",x"c92d7251",x"8ac92d8b",x"8d2d843d",x"0d04fe3d",x"0d800b9e",x"b40c8af8",x"2d818151",x"8ac92d9e",x"84538f52",x"72708105",x"5433518a",x"c92dff12",x"5271ff2e",x"098106ec",x"388b8d2d",x"843d0d04",x"fe3d0d80",x"0b9eb40c",x"8af82d81",x"82518ac9",x"2d80d080",x"8084528b",x"ee2d81f9",x"0a0b80d0",x"80809c0c",x"71087252",x"538bd22d",x"729ebc0c",x"72902a51",x"8ac92d9e",x"bc08882a",x"518ac92d",x"9ebc0851",x"8ac92d8e",x"bf2d8808",x"518ac92d",x"8b8d2d84",x"3d0d0480",x"3d0d810b",x"9eb80c80",x"0b83900a",x"0c85518e",x"aa2d823d",x"0d04803d",x"0d800b9e",x"b80c8bae",x"2d86518e",x"aa2d823d",x"0d04fd3d",x"0d80d080",x"8084548a",x"518eaa2d",x"8bee2d9e",x"a8745253",x"8c942d72",x"88081010",x"80dc8084",x"05717084",x"05530c52",x"fb8084a1",x"ad720c9e",x"840b8814",x"0c73518b",x"d22d8a8e",x"2d8c852d",x"fc3d0d80",x"d0808084",x"7052558b",x"d22d8bee",x"2d8b750c",x"7680d080",x"80940c80",x"750ca080",x"54775383",x"d00a5274",x"518cb42d",x"74518bd2",x"2d8a8e2d",x"8c852dff",x"ab3d0d80",x"0b9eb80c",x"800b9eb4",x"0c800b8e",x"8d0ba080",x"0c5780c4",x"80808455",x"8480b575",x"0c80c880",x"80a453fb",x"ffff7308",x"70720675",x"0c535480",x"c8808094",x"70087076",x"06720c53",x"53a87099",x"85717084",x"05530c99",x"e2710c53",x"9afb0b88",x"120c9c8a",x"0b8c120c",x"93bc0b90",x"120c5388",x"0b80c080",x"80840c90",x"0a538173",x"0c8bae2d",x"fe88880b",x"80dc8080",x"840c81f2",x"0b80d00a",x"0c80d080",x"80847052",x"528bd22d",x"8bee2d71",x"518bd22d",x"76777675",x"933d4141",x"5b5b5b83",x"d00a5c78",x"08708106",x"5152719d",x"389eb808",x"5372f038",x"9eb40852",x"87e87227",x"e638727e",x"0c728390",x"0a0c97a6",x"2d82900a",x"08537980",x"2e81b438",x"7280fe2e",x"09810680",x"f4387680",x"2ec13880",x"7d785856",x"5a827727",x"ffb53883",x"ffff7c0c",x"79fe1853",x"53797227",x"983880dc",x"80808872",x"55587215",x"7033790c",x"52811353",x"737326f2",x"38ff1675",x"11547505",x"ff057033",x"74337072",x"882b077f",x"08535155",x"51527173",x"2e098106",x"feed3874",x"3353728a",x"26fee438",x"7210109d",x"d8057552",x"70085152",x"712dfed3",x"397280fd",x"2e098106",x"8638815b",x"fec53976",x"829f269e",x"387a802e",x"87388073",x"a032545b",x"80d73d77",x"05fde005",x"52727234",x"811757fe",x"a239805a",x"fe9d3972",x"80fe2e09",x"8106fe93",x"387957ff",x"7c0c8177",x"5c5afe87",x"39ff3d0d",x"97dd2d80",x"52805193",x"f32d833d",x"0d049fff",x"fff80d8c",x"ef049fff",x"fff80da0",x"88048808",x"80c08080",x"8808a080",x"082d5088",x"0c810b90",x"0a0c0400",x"00000000",x"820b80c0",x"8080900c",x"0b0b0b04",x"0083f00a",x"0b800ba0",x"80721208",x"720c8412",x"5271712e",x"ff05f238",x"028c050d",x"97d00400",x"00000000",x"00000000",x"00000000",x"00fb3d0d",x"77795555",x"80567575",x"24ab3880",x"74249d38",x"80537352",x"745180e1",x"3f880854",x"75802e85",x"38880830",x"5473880c",x"873d0d04",x"73307681",x"325754dc",x"39743055",x"81567380",x"25d238ec",x"39fa3d0d",x"787a5755",x"80577675",x"24a43875",x"9f2c5481",x"53757432",x"74315274",x"519b3f88",x"08547680",x"2e853888",x"08305473",x"880c883d",x"0d047430",x"558157d7",x"39fc3d0d",x"76785354",x"81538074",x"73265255",x"72802e98",x"3870802e",x"a9388072",x"24a43871",x"10731075",x"72265354",x"5272ea38",x"73517883",x"38745170",x"880c863d",x"0d047281",x"2a72812a",x"53537280",x"2ee63871",x"7426ef38",x"73723175",x"74077481",x"2a74812a",x"55555654",x"e539fc3d",x"0d767079",x"7b555555",x"558f7227",x"8c387275",x"07830651",x"70802ea7",x"38ff1252",x"71ff2e98",x"38727081",x"05543374",x"70810556",x"34ff1252",x"71ff2e09",x"8106ea38",x"74880c86",x"3d0d0474",x"51727084",x"05540871",x"70840553",x"0c727084",x"05540871",x"70840553",x"0c727084",x"05540871",x"70840553",x"0c727084",x"05540871",x"70840553",x"0cf01252",x"718f26c9",x"38837227",x"95387270",x"84055408",x"71708405",x"530cfc12",x"52718326",x"ed387054",x"ff8339fc",x"3d0d7679",x"71028c05",x"9f053357",x"55535583",x"72278a38",x"74830651",x"70802ea2",x"38ff1252",x"71ff2e93",x"38737370",x"81055534",x"ff125271",x"ff2e0981",x"06ef3874",x"880c863d",x"0d047474",x"882b7507",x"7071902b",x"07515451",x"8f7227a5",x"38727170",x"8405530c",x"72717084",x"05530c72",x"71708405",x"530c7271",x"70840553",x"0cf01252",x"718f26dd",x"38837227",x"90387271",x"70840553",x"0cfc1252",x"718326f2",x"387053ff",x"9039fb3d",x"0d777970",x"72078306",x"53545270",x"93387173",x"73085456",x"54717308",x"2e80c438",x"73755452",x"71337081",x"ff065254",x"70802e9d",x"38723355",x"70752e09",x"81069538",x"81128114",x"71337081",x"ff065456",x"545270e5",x"38723355",x"7381ff06",x"7581ff06",x"71713188",x"0c525287",x"3d0d0471",x"0970f7fb",x"fdff1406",x"70f88482",x"81800651",x"51517097",x"38841484",x"16710854",x"56547175",x"082edc38",x"73755452",x"ff963980",x"0b880c87",x"3d0d04ff",x"3d0d9ec4",x"0bfc0570",x"08525270",x"ff2e9138",x"702dfc12",x"70085252",x"70ff2e09",x"8106f138",x"833d0d04",x"04ebe13f",x"04000000",x"00ffffff",x"ff00ffff",x"ffff00ff",x"ffffff00",x"000008c6",x"000008f8",x"000008a0",x"000007b9",x"0000094f",x"00000966",x"0000084c",x"0000084d",x"00000765",x"0000097a",x"01091700",x"00ffef80",x"05f5e100",x"ba011a00",x"00000000",x"00000000",x"00000000",x"00000f4c",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"ffffffff",x"00000000",x"ffffffff",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000");

begin

  process (clk)
  begin
    if rising_edge(clk) then
      if ENA='1' then
        if WEA='1' then
          RAM(conv_integer(ADDRA) ) := DIA;
        end if;
        DOA <= RAM(conv_integer(ADDRA)) ;
      end if;
    end if;
  end process;  

  process (clk)
  begin
    if rising_edge(clk) then
      if ENB='1' then
        if WEB='1' then
          RAM( conv_integer(ADDRB) ) := DIB;
        end if;
        DOB <= RAM(conv_integer(ADDRB)) ;
      end if;
    end if;
  end process;  
end behave;
