library IEEE;
use IEEE.std_logic_1164.all; 
use IEEE.std_logic_unsigned.all; 
use ieee.numeric_std.all;

entity bootloader_dp_32 is
  port (
    CLK:              in std_logic;
    WEA:  in std_logic;
    ENA:  in std_logic;
    MASKA:    in std_logic_vector(3 downto 0);
    ADDRA:         in std_logic_vector(11 downto 2);
    DIA:        in std_logic_vector(31 downto 0);
    DOA:         out std_logic_vector(31 downto 0);
    WEB:  in std_logic;
    ENB:  in std_logic;
    ADDRB:         in std_logic_vector(11 downto 2);
    DIB:        in std_logic_vector(31 downto 0);
    MASKB:    in std_logic_vector(3 downto 0);
    DOB:         out std_logic_vector(31 downto 0)
  );
end entity bootloader_dp_32;

architecture behave of bootloader_dp_32 is

  subtype RAM_WORD is STD_LOGIC_VECTOR (31 downto 0);
  type RAM_TABLE is array (0 to 1023) of RAM_WORD;
 shared variable RAM: RAM_TABLE := RAM_TABLE'(
x"0b0b0b9b",x"c5040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b9b",x"af040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fd0608",x"72830609",x"81058205",x"832b2a83",x"ffff0652",x"04000000",x"00000000",x"00000000",x"71fd0608",x"83ffff73",x"83060981",x"05820583",x"2b2b0906",x"7383ffff",x"0b0b0b0b",x"83a70400",x"72098105",x"72057373",x"09060906",x"73097306",x"070a8106",x"53510400",x"00000000",x"00000000",x"72722473",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71737109",x"71068106",x"30720a10",x"0a720a10",x"0a31050a",x"81065151",x"53510400",x"00000000",x"72722673",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"cc040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"720a722b",x"0a535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72729f06",x"0981050b",x"0b0b88af",x"05040000",x"00000000",x"00000000",x"00000000",x"00000000",x"72722aff",x"739f062a",x"0974090a",x"8106ff05",x"06075351",x"04000000",x"00000000",x"00000000",x"71715351",x"020d0406",x"73830609",x"81058205",x"832b0b2b",x"0772fc06",x"0c515104",x"00000000",x"72098105",x"72050970",x"81050906",x"0a810653",x"51040000",x"00000000",x"00000000",x"00000000",x"72098105",x"72050970",x"81050906",x"0a098106",x"53510400",x"00000000",x"00000000",x"00000000",x"71098105",x"52040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72720981",x"05055351",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097206",x"73730906",x"07535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fc0608",x"72830609",x"81058305",x"1010102a",x"81ff0652",x"04000000",x"00000000",x"00000000",x"71fc0608",x"0b0b0b9e",x"8c738306",x"10100508",x"060b0b0b",x"88b20400",x"00000000",x"00000000",x"0b0b0b89",x"80040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"e8040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097081",x"0509060a",x"8106ff05",x"70547106",x"73097274",x"05ff0506",x"07515151",x"04000000",x"72097081",x"0509060a",x"098106ff",x"05705471",x"06730972",x"7405ff05",x"06075151",x"51040000",x"05ff0504",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"810b0b0b",x"0b9ec80c",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71810552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"02840572",x"10100552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"717105ff",x"05715351",x"020d0400",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"81d53f95",x"e53f0400",x"00000000",x"00000000",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101053",x"51047381",x"ff067383",x"06098105",x"83051010",x"102b0772",x"fc060c51",x"51043c04",x"72728072",x"8106ff05",x"09720605",x"71105272",x"0a100a53",x"72ed3851",x"51535104",x"88088c08",x"90087575",x"9ce42d50",x"50880856",x"900c8c0c",x"880c5104",x"88088c08",x"90087575",x"9ca92d50",x"50880856",x"900c8c0c",x"880c5104",x"88088c08",x"90088eb9",x"2d900c8c",x"0c880c04",x"ff3d0d0b",x"0b80c080",x"3351709e",x"389ed408",x"70085252",x"70802e8a",x"3884129e",x"d40c702d",x"ec39810b",x"0b0b80c0",x"8034833d",x"0d040480",x"3d0d0b0b",x"0b9efc08",x"802e9738",x"0b0b0b0b",x"800b802e",x"8d380b0b",x"0b9efc51",x"0b0b0bf6",x"873f823d",x"0d0404ff",x"3d0d80c4",x"80808452",x"71087082",x"2a708106",x"51515170",x"f338833d",x"0d04ff3d",x"0d80c480",x"80845271",x"0870812a",x"70810651",x"515170f3",x"38738290",x"0a0c833d",x"0d04fe3d",x"0d747080",x"dc808088",x"0c7081ff",x"06ff8311",x"54515371",x"81268d38",x"80fd518a",x"9a2d72a0",x"32518339",x"72518a9a",x"2d843d0d",x"04ff3d0d",x"028f0533",x"5283ffff",x"0b83d00a",x"0c80fe51",x"8a9a2d71",x"518aba2d",x"833d0d04",x"fe3d0d83",x"d00a0870",x"81ff0652",x"528aba2d",x"71882a51",x"8aba2d80",x"fe518a9a",x"2d80c0a0",x"33810587",x"06527180",x"c0a03484",x"3d0d04fe",x"3d0d80c0",x"a4337083",x"2b820781",x"fa065253",x"8ae92d8b",x"882d843d",x"0d04fe3d",x"0d80c0a4",x"3370832b",x"810781f9",x"0652538a",x"e92d8b88",x"2d843d0d",x"0482f6ff",x"0b80cc80",x"80880c80",x"0b80cc80",x"80840c9f",x"0b83900a",x"0c04ff3d",x"0d737008",x"515180c8",x"80808470",x"08708480",x"8007720c",x"5252833d",x"0d04ff3d",x"0d80c880",x"80847008",x"70fbffff",x"06720c52",x"52833d0d",x"04a0900b",x"80ccb40c",x"80c0840b",x"80ccb80c",x"9ba62dff",x"3d0d7351",x"8b710c90",x"11529880",x"80720c80",x"720c7008",x"83ffff06",x"880c833d",x"0d04fa3d",x"0d787a7d",x"ff1e5656",x"585572ff",x"2ea73880",x"56845275",x"750c7408",x"88180cff",x"125271f3",x"38738415",x"7608720c",x"ff155555",x"5272ff2e",x"098106dd",x"38883d0d",x"04f93d0d",x"80d08080",x"845783d0",x"0a588ca2",x"2d76518c",x"cb2d80c0",x"84708808",x"84299880",x"84057170",x"8405530c",x"5656fb80",x"84a1ad75",x"0c9ed80b",x"88170c80",x"70780c77",x"0c760870",x"83ffff06",x"515683ff",x"ff780ca0",x"80548808",x"53775276",x"518cea2d",x"76518c86",x"2d770855",x"75752e89",x"3880c351",x"8a9a2dff",x"39a08408",x"5574fba0",x"90ae802e",x"893880c2",x"518a9a2d",x"ff3980d0",x"0a700870",x"ffbf0672",x"0c565689",x"ff2d8cb9",x"2dff3d0d",x"80c09408",x"811180c0",x"940c5183",x"900a7008",x"70feff06",x"720c5252",x"833d0d04",x"fe3d0d80",x"c0a03370",x"832b8180",x"0780c0a4",x"337181f8",x"06075353",x"538ae92d",x"74818007",x"518aba2d",x"8b882d84",x"3d0d04fe",x"3d0d80d0",x"80808453",x"8ca22d85",x"730c8073",x"0c720870",x"81ff0674",x"5351528c",x"862d7188",x"0c843d0d",x"04fc3d0d",x"76811133",x"82123371",x"81800a29",x"71848080",x"29058314",x"33708280",x"29128416",x"33527105",x"a0800586",x"16851733",x"57525353",x"55575553",x"ff135372",x"ff2e9138",x"73708105",x"55335271",x"75708105",x"5734e939",x"89518ed8",x"2d863d0d",x"04f93d0d",x"795680d0",x"80808457",x"8ca22d81",x"16338217",x"33718280",x"29055353",x"71802e94",x"38851672",x"55537270",x"81055433",x"770cff14",x"5473f338",x"83163384",x"17337182",x"80290556",x"52805473",x"75279738",x"73587777",x"0c731677",x"08535371",x"73348114",x"54747426",x"ed387651",x"8c862d80",x"c0a03370",x"832b8180",x"0780c0a4",x"337181f8",x"06075353",x"548ae92d",x"8184518a",x"ba2d7488",x"2a518aba",x"2d74518a",x"ba2d8054",x"7375278f",x"38731670",x"3352528a",x"ba2d8114",x"54ee398b",x"882d893d",x"0d04fc3d",x"0d80d080",x"80840b81",x"1854558b",x"b72d8ca2",x"2d86750c",x"74518c86",x"2d8ca22d",x"82750c72",x"70810554",x"33750c72",x"70810554",x"33750c72",x"70810554",x"33750c81",x"ff547270",x"81055433",x"750cff14",x"54738025",x"f1387451",x"8c862d8f",x"832d8808",x"81065271",x"f638863d",x"0d04fa3d",x"0d785680",x"d0808084",x"548ca22d",x"86740c73",x"518c862d",x"8ca22d81",x"ad740c81",x"16338217",x"33718280",x"29058318",x"33760c84",x"1833760c",x"85183376",x"0c585280",x"55747727",x"af387480",x"2e88388c",x"a22d81ad",x"740c7416",x"86113375",x"0c871133",x"750c5273",x"518c862d",x"8f832d88",x"08810652",x"71f63882",x"1555ce39",x"8ca22d84",x"740c7351",x"8c862d80",x"c0a03370",x"832b8180",x"0780c0a4",x"337181f8",x"06075353",x"538ae92d",x"8187518a",x"ba2d8b88",x"2d883d0d",x"04fc3d0d",x"76811133",x"82123371",x"902b7188",x"2b078314",x"33707207",x"882b8416",x"33710751",x"52535657",x"55528851",x"8ed82d81",x"ff518a9a",x"2d80c480",x"80845473",x"0870812a",x"70810651",x"515271f3",x"38728480",x"800780c4",x"8080840c",x"863d0d04",x"fd3d0d8f",x"832d8808",x"88088106",x"535371f3",x"3880c0a0",x"3370832b",x"81800780",x"c0a43371",x"81f80607",x"5353548a",x"e92d8183",x"518aba2d",x"72518aba",x"2d8b882d",x"853d0d04",x"fe3d0d80",x"0b80c094",x"0c80c0a0",x"3370832b",x"81800780",x"c0a43371",x"81f80607",x"5353538a",x"e92d8181",x"518aba2d",x"9ed85393",x"52727081",x"05543351",x"8aba2dff",x"125271ff",x"2e098106",x"ec388b88",x"2d843d0d",x"04fe3d0d",x"800b80c0",x"940c80c0",x"a0337083",x"2b818007",x"80c0a433",x"7181f806",x"07535353",x"8ae92d81",x"82518aba",x"2d80d080",x"8084528c",x"a22d81f9",x"0a0b80d0",x"80809c0c",x"71087252",x"538c862d",x"7280c0a8",x"0c72902a",x"518aba2d",x"80c0a808",x"882a518a",x"ba2d80c0",x"a808518a",x"ba2d8f83",x"2d880851",x"8aba2d8b",x"882d843d",x"0d04803d",x"0d810b80",x"c0980c80",x"0b83900a",x"0c85518e",x"d82d823d",x"0d04803d",x"0d800b80",x"c0980c8b",x"ed2d8651",x"8ed82d82",x"3d0d04fd",x"3d0d80d0",x"80808454",x"8a518ed8",x"2d8ca22d",x"80c08474",x"52538ccb",x"2d728808",x"84299880",x"84057170",x"8405530c",x"52fb8084",x"a1ad720c",x"9ed80b88",x"140c7351",x"8c862d89",x"ff2d8cb9",x"2dffb13d",x"0d80d33d",x"0856800b",x"80c0980c",x"800b80c0",x"940c800b",x"df80179e",x"dd71902a",x"71565657",x"55577272",x"70810554",x"3473882a",x"53727234",x"73821634",x"75982a52",x"718b1634",x"75902a52",x"718c1634",x"75882a52",x"718d1634",x"758e1634",x"7680c090",x"348eb90b",x"80ccb40c",x"8480b30b",x"80c48080",x"840c80c8",x"8080a453",x"fbffff73",x"08707206",x"750c5354",x"80c88080",x"94700870",x"7606720c",x"5353880b",x"80c08080",x"840c810b",x"900a0c8b",x"ed2dfe88",x"880b80dc",x"8080840c",x"81f20b80",x"d00a0c80",x"d0808084",x"7052528c",x"862d8ca2",x"2d71518c",x"862d8ca2",x"2d84720c",x"71518c86",x"2d767757",x"5580c480",x"80840870",x"81065152",x"71a03880",x"c0980853",x"72eb3880",x"c0940852",x"87e87227",x"e0387290",x"0a0c7283",x"900a0c9b",x"9e2d8290",x"0a085375",x"802e8294",x"387280fe",x"2e098106",x"81cd3876",x"802effb9",x"38800b8a",x"3d555682",x"7727ffad",x"3883d00a",x"08527176",x"2e87388b",x"d22dff9d",x"39733370",x"872a8132",x"53537180",x"2e993872",x"87065271",x"ff873875",x"80c0a434",x"7580c0a0",x"348bb72d",x"fef73972",x"b8067083",x"2a80c0a4",x"33555152",x"71732e80",x"c0388bd2",x"2d80c0a4",x"3380c09c",x"3480c0a4",x"33720587",x"06708281",x"2980c0ac",x"05ff1955",x"515272ff",x"2e923873",x"70810555",x"33727081",x"055434ff",x"1353eb39",x"810b80c0",x"9034fea5",x"39811387",x"06527180",x"c0a43475",x"80c09033",x"53537183",x"38735381",x"13335271",x"8b26fe85",x"38718429",x"9e980581",x"14527008",x"5152712d",x"fdf33972",x"80fd2e09",x"81068638",x"8155fde5",x"3976829f",x"26a53874",x"802e8738",x"8073a032",x"54557280",x"dc808088",x"0c80d13d",x"7705fde0",x"05527272",x"34811757",x"fdbb3980",x"56fdb639",x"7280fe2e",x"098106fd",x"ac387557",x"ff0b83d0",x"0a0c8177",x"5656fd9d",x"39ff3d0d",x"9bfd2d73",x"52805196",x"dd2d833d",x"0d0483ff",x"fff80d8d",x"a50483ff",x"fff80d80",x"ccbc0488",x"0880c080",x"80880880",x"ccb4082d",x"50880c81",x"0b900a0c",x"0480700c",x"faad95b4",x"da0b8180",x"8071710c",x"7180082e",x"87387011",x"519bd104",x"519b8d2d",x"00000000",x"00000000",x"00000000",x"820b80c0",x"8080900c",x"0b0b0b04",x"0083f00a",x"0b800ba0",x"80721208",x"720c8412",x"5271712e",x"ff05f238",x"028c050d",x"9bf00400",x"00000000",x"00000000",x"00000000",x"00fb3d0d",x"77795555",x"80567476",x"25863874",x"30558156",x"73802588",x"38733076",x"81325754",x"80537352",x"745180ca",x"3f880854",x"75802e85",x"38880830",x"5473880c",x"873d0d04",x"fa3d0d78",x"7a575580",x"57747725",x"86387430",x"55815775",x"9f2c5481",x"53757432",x"74315274",x"51943f88",x"08547680",x"2e853888",x"08305473",x"880c883d",x"0d04fc3d",x"0d767853",x"54815380",x"55873971",x"10731054",x"52737226",x"5172802e",x"a7387080",x"2e863871",x"8025e838",x"72802e98",x"38717426",x"89387372",x"31757407",x"56547281",x"2a72812a",x"5353e539",x"73517883",x"38745170",x"880c863d",x"0d04ff3d",x"0d9ef00b",x"fc055271",x"08ff2e8b",x"38710851",x"702dfc12",x"52f13983",x"3d0d0404",x"eb9e3f04",x"00ffffff",x"ff00ffff",x"ffff00ff",x"ffffff00",x"00000a34",x"00000a7d",x"000009f8",x"000007fd",x"00000aee",x"00000b06",x"00000906",x"000009a5",x"000007a9",x"00000b1b",x"000008a6",x"00000000",x"00000000",x"00000000",x"00000f78",x"01090600",x"00000000",x"05b8d800",x"b4041700",x"00000000",x"ffffffff",x"00000000",x"ffffffff",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000");

begin

  process (clk)
  begin
    if rising_edge(clk) then
      if ENA='1' then
        if WEA='1' then
          RAM(conv_integer(ADDRA) ) := DIA;
        end if;
        DOA <= RAM(conv_integer(ADDRA)) ;
      end if;
    end if;
  end process;  

  process (clk)
  begin
    if rising_edge(clk) then
      if ENB='1' then
        if WEB='1' then
          RAM( conv_integer(ADDRB) ) := DIB;
        end if;
        DOB <= RAM(conv_integer(ADDRB)) ;
      end if;
    end if;
  end process;  
end behave;
