library IEEE;
use IEEE.std_logic_1164.all; 
use IEEE.std_logic_unsigned.all; 
use ieee.numeric_std.all;

entity bootloader_dp_32 is
  port (
    CLK:              in std_logic;
    WEA:  in std_logic;
    ENA:  in std_logic;
    MASKA:    in std_logic_vector(3 downto 0);
    ADDRA:         in std_logic_vector(11 downto 2);
    DIA:        in std_logic_vector(31 downto 0);
    DOA:         out std_logic_vector(31 downto 0);
    WEB:  in std_logic;
    ENB:  in std_logic;
    ADDRB:         in std_logic_vector(11 downto 2);
    DIB:        in std_logic_vector(31 downto 0);
    MASKB:    in std_logic_vector(3 downto 0);
    DOB:         out std_logic_vector(31 downto 0)
  );
end entity bootloader_dp_32;

architecture behave of bootloader_dp_32 is

  subtype RAM_WORD is STD_LOGIC_VECTOR (31 downto 0);
  type RAM_TABLE is array (0 to 1023) of RAM_WORD;
 shared variable RAM: RAM_TABLE := RAM_TABLE'(
x"0b0b0b98",x"9b040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b98",x"86040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fd0608",x"72830609",x"81058205",x"832b2a83",x"ffff0652",x"04000000",x"00000000",x"00000000",x"71fd0608",x"83ffff73",x"83060981",x"05820583",x"2b2b0906",x"7383ffff",x"0b0b0b0b",x"83a70400",x"72098105",x"72057373",x"09060906",x"73097306",x"070a8106",x"53510400",x"00000000",x"00000000",x"72722473",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71737109",x"71068106",x"30720a10",x"0a720a10",x"0a31050a",x"81065151",x"53510400",x"00000000",x"72722673",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"cc040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"720a722b",x"0a535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72729f06",x"0981050b",x"0b0b88af",x"05040000",x"00000000",x"00000000",x"00000000",x"00000000",x"72722aff",x"739f062a",x"0974090a",x"8106ff05",x"06075351",x"04000000",x"00000000",x"00000000",x"71715351",x"020d0406",x"73830609",x"81058205",x"832b0b2b",x"0772fc06",x"0c515104",x"00000000",x"72098105",x"72050970",x"81050906",x"0a810653",x"51040000",x"00000000",x"00000000",x"00000000",x"72098105",x"72050970",x"81050906",x"0a098106",x"53510400",x"00000000",x"00000000",x"00000000",x"71098105",x"52040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72720981",x"05055351",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097206",x"73730906",x"07535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fc0608",x"72830609",x"81058305",x"1010102a",x"81ff0652",x"04000000",x"00000000",x"00000000",x"71fc0608",x"0b0b0b9a",x"fc738306",x"10100508",x"060b0b0b",x"88b20400",x"00000000",x"00000000",x"0b0b0b89",x"80040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"e8040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097081",x"0509060a",x"8106ff05",x"70547106",x"73097274",x"05ff0506",x"07515151",x"04000000",x"72097081",x"0509060a",x"098106ff",x"05705471",x"06730972",x"7405ff05",x"06075151",x"51040000",x"05ff0504",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"810b0b0b",x"0b9bb40c",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71810552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"02840572",x"10100552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"717105ff",x"05715351",x"020d0400",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"81dd3f92",x"cd3f0400",x"00000000",x"00000000",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101053",x"51047381",x"ff067383",x"06098105",x"83051010",x"102b0772",x"fc060c51",x"51043c04",x"72728072",x"8106ff05",x"09720605",x"71105272",x"0a100a53",x"72ed3851",x"51535104",x"88088c08",x"90087575",x"99bd2d50",x"50880856",x"900c8c0c",x"880c5104",x"88088c08",x"90087575",x"98f92d50",x"50880856",x"900c8c0c",x"880c5104",x"88088c08",x"90088df6",x"2d900c8c",x"0c880c04",x"ff3d0d0b",x"0b0b9bd8",x"335170a6",x"389bc008",x"70085252",x"70802e92",x"3884129b",x"c00c702d",x"9bc00870",x"08525270",x"f038810b",x"0b0b0b9b",x"d834833d",x"0d040480",x"3d0d0b0b",x"0b9c8408",x"802e8e38",x"0b0b0b0b",x"800b802e",x"09810685",x"38823d0d",x"040b0b0b",x"9c84510b",x"0b0bf5f8",x"3f823d0d",x"0404ff3d",x"0d80c480",x"80845271",x"0870822a",x"70810651",x"515170f3",x"38833d0d",x"04ff3d0d",x"80c48080",x"84527108",x"70812a70",x"81065151",x"5170f338",x"7382900a",x"0c833d0d",x"04fe3d0d",x"747080dc",x"8080880c",x"7081ff06",x"ff831154",x"51537181",x"268d3880",x"fd518aa9",x"2d72a032",x"51833972",x"518aa92d",x"843d0d04",x"803d0d83",x"ffff0b83",x"d00a0c80",x"fe518aa9",x"2d823d0d",x"04ff3d0d",x"83d00a08",x"70882a52",x"528ac92d",x"7181ff06",x"518ac92d",x"80fe518a",x"a92d833d",x"0d0482f6",x"ff0b80cc",x"8080880c",x"800b80cc",x"8080840c",x"9f0b8390",x"0a0c04ff",x"3d0d7370",x"08515180",x"c8808084",x"70087084",x"80800772",x"0c525283",x"3d0d04ff",x"3d0d80c8",x"80808470",x"0870fbff",x"ff06720c",x"5252833d",x"0d04a090",x"0ba0800c",x"9bdc0ba0",x"840c97fe",x"2dff3d0d",x"73518b71",x"0c901152",x"98808072",x"0c80720c",x"700883ff",x"ff06880c",x"833d0d04",x"fa3d0d78",x"7a7dff1e",x"57575853",x"73ff2ea7",x"38805684",x"5275730c",x"72088818",x"0cff1252",x"71f33874",x"84167408",x"720cff16",x"56565273",x"ff2e0981",x"06dd3888",x"3d0d04f9",x"3d0d80d0",x"80808456",x"83d00a58",x"8be32d75",x"518c892d",x"9bdc7088",x"08101098",x"80840571",x"70840553",x"0c5657fb",x"8084a1ad",x"750c9bc4",x"0b88180c",x"8070770c",x"760c7508",x"7083ffff",x"06515783",x"ffff780c",x"a0805488",x"08537752",x"75518ca8",x"2d75518b",x"c72d7708",x"5574772e",x"893880c3",x"518aa92d",x"ff39a084",x"085574fb",x"a08cae80",x"2e893880",x"c2518aa9",x"2dff3980",x"d00a7008",x"70ffbf06",x"720c5656",x"8a8e2d8b",x"fa2dff3d",x"0d9be808",x"81119be8",x"0c518390",x"0a700870",x"feff0672",x"0c525283",x"3d0d0480",x"3d0d8af8",x"2d728180",x"07518ac9",x"2d8b8d2d",x"823d0d04",x"fe3d0d80",x"d0808084",x"538be32d",x"85730c80",x"730c7208",x"7081ff06",x"74535152",x"8bc72d71",x"880c843d",x"0d04fc3d",x"0d768111",x"33821233",x"7181800a",x"29718480",x"80290583",x"14337082",x"80291284",x"16335271",x"05a08005",x"86168517",x"33575253",x"53555755",x"53ff1353",x"72ff2e91",x"38737081",x"05553352",x"71757081",x"055734e9",x"3989518e",x"932d863d",x"0d04f93d",x"0d795780",x"d0808084",x"568be32d",x"81173382",x"18337182",x"80290553",x"5371802e",x"94388517",x"72555372",x"70810554",x"33760cff",x"145473f3",x"38831733",x"84183371",x"82802905",x"56528054",x"73752797",x"38735877",x"760c7317",x"76085353",x"71733481",x"14547474",x"26ed3875",x"518bc72d",x"8af82d81",x"84518ac9",x"2d74882a",x"518ac92d",x"74518ac9",x"2d805473",x"75278f38",x"73177033",x"52528ac9",x"2d811454",x"ee398b8d",x"2d893d0d",x"04f93d0d",x"795680d0",x"80808455",x"8be32d86",x"750c7451",x"8bc72d8b",x"e32d81ad",x"70760c81",x"17338218",x"33718280",x"29058319",x"33780c84",x"1933780c",x"85193378",x"0c595353",x"80547377",x"27b33872",x"5873802e",x"87388be3",x"2d77750c",x"73168611",x"33760c87",x"1133760c",x"5274518b",x"c72d8ea8",x"2d880881",x"065271f6",x"38821454",x"767426d1",x"388be32d",x"84750c74",x"518bc72d",x"8af82d81",x"87518ac9",x"2d8b8d2d",x"893d0d04",x"fc3d0d76",x"81113382",x"12337190",x"2b71882b",x"07831433",x"70720788",x"2b841633",x"71075152",x"53575754",x"5288518e",x"932d81ff",x"518aa92d",x"80c48080",x"84537208",x"70812a70",x"81065151",x"5271f338",x"73848080",x"0780c480",x"80840c86",x"3d0d04fe",x"3d0d8ea8",x"2d880888",x"08810653",x"5371f338",x"8af82d81",x"83518ac9",x"2d72518a",x"c92d8b8d",x"2d843d0d",x"04fe3d0d",x"800b9be8",x"0c8af82d",x"8181518a",x"c92d9bc4",x"53935272",x"70810554",x"33518ac9",x"2dff1252",x"71ff2e09",x"8106ec38",x"8b8d2d84",x"3d0d04fe",x"3d0d800b",x"9be80c8a",x"f82d8182",x"518ac92d",x"80d08080",x"84528be3",x"2d81f90a",x"0b80d080",x"809c0c71",x"08725253",x"8bc72d72",x"9bf00c72",x"902a518a",x"c92d9bf0",x"08882a51",x"8ac92d9b",x"f008518a",x"c92d8ea8",x"2d880851",x"8ac92d8b",x"8d2d843d",x"0d04803d",x"0d810b9b",x"ec0c800b",x"83900a0c",x"85518e93",x"2d823d0d",x"04803d0d",x"800b9bec",x"0c8bae2d",x"86518e93",x"2d823d0d",x"04fd3d0d",x"80d08080",x"84548a51",x"8e932d8b",x"e32d9bdc",x"7452538c",x"892d7288",x"08101098",x"80840571",x"70840553",x"0c52fb80",x"84a1ad72",x"0c9bc40b",x"88140c73",x"518bc72d",x"8a8e2d8b",x"fa2dffab",x"3d0d80d9",x"3d085680",x"0b9bec0c",x"800b9be8",x"0c800bdf",x"80179bc9",x"71902a71",x"56565755",x"57727270",x"81055434",x"73882a53",x"72723473",x"82163475",x"8b16348d",x"f60ba080",x"0c80c480",x"80845584",x"80b3750c",x"80c88080",x"a453fbff",x"ff730870",x"7206750c",x"535480c8",x"80809470",x"08707606",x"720c5353",x"880b80c0",x"8080840c",x"900a5381",x"730c8bae",x"2dfe8888",x"0b80dc80",x"80840c81",x"f20b80d0",x"0a0c80d0",x"80808470",x"52528bc7",x"2d8be32d",x"71518bc7",x"2d8be32d",x"84720c71",x"518bc72d",x"76777675",x"933d4141",x"5b5b5b83",x"d00a5c78",x"08708106",x"5152719d",x"389bec08",x"5372f038",x"9be80852",x"87e87227",x"e638727e",x"0c728390",x"0a0c97f6",x"2d82900a",x"08537980",x"2e81b438",x"7280fe2e",x"09810680",x"f4387680",x"2ec13880",x"7d785757",x"5a827727",x"ffb53883",x"ffff7c0c",x"79fe1853",x"53797227",x"983880dc",x"80808872",x"55587216",x"7033790c",x"52811353",x"737326f2",x"38ff1576",x"11547605",x"ff057033",x"74337072",x"882b077f",x"08535155",x"51527173",x"2e098106",x"feed3875",x"3353728a",x"26fee438",x"7210109b",x"88057652",x"70085152",x"712dfed3",x"397280fd",x"2e098106",x"8638815b",x"fec53976",x"829f269e",x"387a802e",x"87388073",x"a032545b",x"80d73d77",x"05fde005",x"52727234",x"811757fe",x"a239805a",x"fe9d3972",x"80fe2e09",x"8106fe93",x"387957ff",x"7c0c8177",x"5c5afe87",x"39ff3d0d",x"98cd2d73",x"52805194",x"b22d833d",x"0d0483ff",x"fff80d8c",x"e30483ff",x"fff80da0",x"88048808",x"80c08080",x"8808a080",x"082d5088",x"0c810b90",x"0a0c0480",x"700cfaad",x"95b4da0b",x"81808071",x"710c7180",x"082e8738",x"70115198",x"a7045197",x"e52d0000",x"00000000",x"820b80c0",x"8080900c",x"0b0b0b04",x"0083f00a",x"0b800ba0",x"80721208",x"720c8412",x"5271712e",x"ff05f238",x"028c050d",x"98c00400",x"00000000",x"00000000",x"00000000",x"00fb3d0d",x"77795555",x"80567575",x"24ab3880",x"74249d38",x"80537352",x"745180e1",x"3f880854",x"75802e85",x"38880830",x"5473880c",x"873d0d04",x"73307681",x"325754dc",x"39743055",x"81567380",x"25d238ec",x"39fa3d0d",x"787a5755",x"80577675",x"24a43875",x"9f2c5481",x"53757432",x"74315274",x"519b3f88",x"08547680",x"2e853888",x"08305473",x"880c883d",x"0d047430",x"558157d7",x"39fc3d0d",x"76785354",x"81538074",x"73265255",x"72802e98",x"3870802e",x"a9388072",x"24a43871",x"10731075",x"72265354",x"5272ea38",x"73517883",x"38745170",x"880c863d",x"0d047281",x"2a72812a",x"53537280",x"2ee63871",x"7426ef38",x"73723175",x"74077481",x"2a74812a",x"55555654",x"e539ff3d",x"0d9bf80b",x"fc057008",x"525270ff",x"2e913870",x"2dfc1270",x"08525270",x"ff2e0981",x"06f13883",x"3d0d0404",x"eeae3f04",x"00ffffff",x"ff00ffff",x"ffff00ff",x"ffffff00",x"0000093d",x"0000096f",x"00000917",x"000007a2",x"000009c6",x"000009dd",x"00000835",x"000008c4",x"0000074e",x"000009f1",x"00000000",x"00000000",x"00000000",x"00000e00",x"01090600",x"00000000",x"05b8d800",x"b4031700",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"ffffffff",x"00000000",x"ffffffff",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000");

begin

  process (clk)
  begin
    if rising_edge(clk) then
      if ENA='1' then
        if WEA='1' then
          RAM(conv_integer(ADDRA) ) := DIA;
        end if;
        DOA <= RAM(conv_integer(ADDRA)) ;
      end if;
    end if;
  end process;  

  process (clk)
  begin
    if rising_edge(clk) then
      if ENB='1' then
        if WEB='1' then
          RAM( conv_integer(ADDRB) ) := DIB;
        end if;
        DOB <= RAM(conv_integer(ADDRB)) ;
      end if;
    end if;
  end process;  
end behave;
