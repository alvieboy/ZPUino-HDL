library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

library work;
use work.zpu_config.all;
use work.zpupkg.all;
use work.zpuinopkg.all;
use work.zpuino_config.all;
use work.wishbonepkg.all;

entity wb_rom_ram is
  port (
    ram_wb_clk_i:       in std_logic;
    ram_wb_rst_i:       in std_logic;
    ram_wb_ack_o:       out std_logic;
    ram_wb_dat_i:       in std_logic_vector(wordSize-1 downto 0);
    ram_wb_dat_o:       out std_logic_vector(wordSize-1 downto 0);
    ram_wb_adr_i:       in std_logic_vector(maxAddrBitIncIO downto 0);
    ram_wb_cyc_i:       in std_logic;
    ram_wb_stb_i:       in std_logic;
    ram_wb_we_i:        in std_logic;

    rom_wb_clk_i:       in std_logic;
    rom_wb_rst_i:       in std_logic;
    rom_wb_ack_o:       out std_logic;
    rom_wb_dat_o:       out std_logic_vector(wordSize-1 downto 0);
    rom_wb_adr_i:       in std_logic_vector(maxAddrBitIncIO downto 0);
    rom_wb_cyc_i:       in std_logic;
    rom_wb_cti_i:       in std_logic_vector(2 downto 0);
    rom_wb_stb_i:       in std_logic;
    rom_wb_stall_o:     out std_logic
  );
end entity wb_rom_ram;


architecture behave of wb_rom_ram is

  component zpuino_icache is
  port (
    wb_clk_i:       in std_logic;
    wb_rst_i:       in std_logic;

    wb_ack_o:       out std_logic;
    wb_dat_o:       out std_logic_vector(wordSize-1 downto 0);
    wb_adr_i:       in std_logic_vector(maxAddrBitIncIO downto 0);
    wb_cyc_i:       in std_logic;
    wb_stb_i:       in std_logic;
    wb_stall_o:     out std_logic;

    -- Master wishbone interface

    m_wb_ack_i:       in std_logic;
    m_wb_dat_i:       in std_logic_vector(wordSize-1 downto 0);
    m_wb_dat_o:       out std_logic_vector(wordSize-1 downto 0);
    m_wb_adr_o:       out std_logic_vector(maxAddrBitIncIO downto 0);
    m_wb_cyc_o:       out std_logic;
    m_wb_stb_o:       out std_logic;
    m_wb_stall_i:     in std_logic;
    m_wb_we_o:        out std_logic
  );
  end component zpuino_icache;

  component dualport_ram is
  generic (
    maxbit: integer
  );
  port (
    clk:              in std_logic;
    memAWriteEnable:  in std_logic;
    memAWriteMask:    in std_logic_vector(3 downto 0);
    memAAddr:         in std_logic_vector(maxbit downto 2);
    memAWrite:        in std_logic_vector(31 downto 0);
    memARead:         out std_logic_vector(31 downto 0);
    memAEnable:       in std_logic;
    memBWriteEnable:  in std_logic;
    memBWriteMask:    in std_logic_vector(3 downto 0);
    memBAddr:         in std_logic_vector(maxbit downto 2);
    memBWrite:        in std_logic_vector(31 downto 0);
    memBRead:         out std_logic_vector(31 downto 0);
    memBEnable:       in std_logic;
    memErr:           out std_logic
  );
  end component dualport_ram;

  constant i_maxAddrBit: integer := 13; -- maxAddrBit


  signal memAWriteEnable:  std_logic;
  signal memAWriteMask:    std_logic_vector(3 downto 0);
  signal memAAddr:         std_logic_vector(i_maxAddrBit downto 2);
  signal memAWrite:        std_logic_vector(31 downto 0);
  signal memARead:         std_logic_vector(31 downto 0);
  signal memAEnable:       std_logic;
  signal memBWriteEnable:  std_logic;
  signal memBWriteMask:    std_logic_vector(3 downto 0);
  signal memBAddr:         std_logic_vector(i_maxAddrBit downto 2);
  signal memBWrite:        std_logic_vector(31 downto 0);
  signal memBRead:         std_logic_vector(31 downto 0);
  signal memBEnable:       std_logic;

  --signal rom_burst: std_logic;
  signal rom_do_wait: std_logic;

  type ramregs_type is record
    do_wait: std_logic;
  end record;
  signal ramregs: ramregs_type;

  signal i_rom_wb_clk_i:       std_logic;
  signal i_rom_wb_rst_i:       std_logic;
  signal i_rom_wb_ack_o:       std_logic;
  signal i_rom_wb_dat_o:       std_logic_vector(wordSize-1 downto 0);
  signal i_rom_wb_adr_i:       std_logic_vector(maxAddrBitIncIO downto 0);
  signal i_rom_wb_cyc_i:       std_logic;
  signal i_rom_wb_stb_i:       std_logic;
  signal i_rom_wb_stall_o:       std_logic;

begin

  -- System ROM/RAM

  ramrom: dualport_ram
  generic map (
    maxbit => 13 --maxAddrBit
  )
  port map (
    clk               => ram_wb_clk_i,
    memAWriteEnable   => memAWriteEnable,
    memAWriteMask     => memAWriteMask,
    memAAddr          => memAAddr,
    memAWrite         => memAWrite,
    memARead          => memARead,
    memAEnable        => memAEnable,
    memBWriteEnable   => memBWriteEnable,
    memBWriteMask     => memBWriteMask,
    memBAddr          => memBAddr,
    memBWrite         => memBWrite,
    memBRead          => memBRead,
    memBEnable        => memBEnable
  );

  memBWrite       <= (others => DontCareValue);
  memBWriteMask   <= (others => DontCareValue);
  memBWriteEnable <= '0';

  i_rom_wb_dat_o    <= memBRead;
  memBAddr        <= i_rom_wb_adr_i(i_maxAddrBit downto 2);
  memBEnable      <= i_rom_wb_cyc_i and i_rom_wb_stb_i;

  icache: zpuino_icache
  port map (
    wb_clk_i    => rom_wb_clk_i,
    wb_rst_i    => rom_wb_rst_i,

    wb_ack_o    => rom_wb_ack_o,
    wb_dat_o    => rom_wb_dat_o,
    wb_adr_i    => rom_wb_adr_i,
    wb_cyc_i    => rom_wb_cyc_i,
    wb_stb_i    => rom_wb_stb_i,
    wb_stall_o  => rom_wb_stall_o,

    -- Master wishbone interface

    m_wb_ack_i  => i_rom_wb_ack_o,
    m_wb_dat_i  => i_rom_wb_dat_o,
    --m_wb_dat_o  => i_rom_wb_dat_i,
    m_wb_adr_o  => i_rom_wb_adr_i,
    m_wb_cyc_o  => i_rom_wb_cyc_i,
    m_wb_stb_o  => i_rom_wb_stb_i,
    --m_wb_we_o   => i_rom_wb_we_i,
    m_wb_stall_i => '0'
  );







  -- ROM ack

  process(rom_wb_clk_i)
  begin
    if rising_edge(rom_wb_clk_i) then
      if rom_wb_rst_i='1' then
        i_rom_wb_ack_o <= '0';
        --rom_burst <= '0';
        rom_do_wait<='0';
      else
        if rom_do_wait='1' then
          if rom_wb_cti_i=CTI_CYCLE_INCRADDR then
              --rom_burst<='1';
              rom_do_wait<='0';
              i_rom_wb_ack_o<='1';
            else
            
              i_rom_wb_ack_o<='0';
              rom_do_wait<='0';
          end if;
        else

          if i_rom_wb_cyc_i='1' and i_rom_wb_stb_i='1' then
            if rom_wb_cti_i=CTI_CYCLE_INCRADDR then
              --rom_burst<='1';
              rom_do_wait<='0';
              i_rom_wb_ack_o<='1';
            else
              --rom_burst<='0';
              rom_do_wait<='1';
              i_rom_wb_ack_o<='1';
            end if;
          elsif i_rom_wb_cyc_i='0' then
            i_rom_wb_ack_o<='0';
          end if;
        end if;
      end if;
    end if;
  end process;

  -- RAM

  memAWrite       <= ram_wb_dat_i;
  memAWriteMask   <= (others => '1');

  ram_wb_dat_o    <= memARead;
  memAAddr        <= ram_wb_adr_i(i_maxAddrBit downto 2);
  memAEnable      <= ram_wb_cyc_i and ram_wb_stb_i;

  -- RAM ack

  process(ram_wb_clk_i, ramregs, ram_wb_rst_i,
          ram_wb_stb_i, ram_wb_cyc_i, ram_wb_we_i)
    variable w: ramregs_type;
  begin

    w:=ramregs;
    --ram_wb_ack_o<='0';
    --memAWriteEnable <= '0';


      ram_wb_ack_o<='0';
      memAWriteEnable <= '0';

      if ramregs.do_wait='1' then
        w.do_wait:='0';
        ram_wb_ack_o<='1';
        if ram_wb_we_i='1' then
          memAWriteEnable <= '1';
        end if;
      else

      if ram_wb_stb_i='1' and ram_wb_cyc_i='1' then
--        if ram_wb_we_i='1' then
--          memAWriteEnable <= '1';
--          ram_wb_ack_o<='1';
--        else
          w.do_wait:='1';
--        end if;
      end if;
      end if;

    if ram_wb_rst_i='1' then
      w.do_wait:='0';
    end if;

    if rising_edge(ram_wb_clk_i) then
      ramregs<=w;
    end if;

  end process;
  
  --ram_wb_ack_o <= '1' when ram_wb_cyc_i='1' and ram_wb_stb_i='1' and ram_wb_we_i='1' else ram_wb_ack_o_i;

end behave;

