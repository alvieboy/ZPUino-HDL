library IEEE;
use IEEE.std_logic_1164.all; 
use IEEE.std_logic_unsigned.all; 
use ieee.numeric_std.all;

entity dualport_ram is
  port (
    clk:              in std_logic;
    memAWriteEnable:  in std_logic;
    memAAddr:         in std_logic_vector(14 downto 2);
    memAWrite:        in std_logic_vector(31 downto 0);
    memARead:         out std_logic_vector(31 downto 0);
    memBWriteEnable:  in std_logic;
    memBAddr:         in std_logic_vector(14 downto 2);
    memBWrite:        in std_logic_vector(31 downto 0);
    memBRead:         out std_logic_vector(31 downto 0)
  );
end entity dualport_ram;

architecture behave of dualport_ram is


  subtype RAM_WORD is STD_LOGIC_VECTOR (31 downto 0);
  type RAM_TABLE is array (0 to 8191) of RAM_WORD;

  shared variable RAM: RAM_TABLE := RAM_TABLE'(
RAM_WORD'(x"0b0b0bb6"),
RAM_WORD'(x"d0700b0b"),
RAM_WORD'(x"8180940c"),
RAM_WORD'(x"3a0b0b0b"),
RAM_WORD'(x"99a00400"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"0b0b0b89"),
RAM_WORD'(x"ab040000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"71fd0608"),
RAM_WORD'(x"72830609"),
RAM_WORD'(x"81058205"),
RAM_WORD'(x"832b2a83"),
RAM_WORD'(x"ffff0652"),
RAM_WORD'(x"04000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"71fd0608"),
RAM_WORD'(x"83ffff73"),
RAM_WORD'(x"83060981"),
RAM_WORD'(x"05820583"),
RAM_WORD'(x"2b2b0906"),
RAM_WORD'(x"7383ffff"),
RAM_WORD'(x"0b0b0b0b"),
RAM_WORD'(x"83a50400"),
RAM_WORD'(x"72098105"),
RAM_WORD'(x"72057373"),
RAM_WORD'(x"09060906"),
RAM_WORD'(x"73097306"),
RAM_WORD'(x"070a8106"),
RAM_WORD'(x"53510400"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"72722473"),
RAM_WORD'(x"732e0753"),
RAM_WORD'(x"51040000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"71737109"),
RAM_WORD'(x"71068106"),
RAM_WORD'(x"30720a10"),
RAM_WORD'(x"0a720a10"),
RAM_WORD'(x"0a31050a"),
RAM_WORD'(x"81065151"),
RAM_WORD'(x"53510400"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"72722673"),
RAM_WORD'(x"732e0753"),
RAM_WORD'(x"51040000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"0b0b0b88"),
RAM_WORD'(x"c3040000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"720a722b"),
RAM_WORD'(x"0a535104"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"72729f06"),
RAM_WORD'(x"0981050b"),
RAM_WORD'(x"0b0b88a6"),
RAM_WORD'(x"05040000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"72722aff"),
RAM_WORD'(x"739f062a"),
RAM_WORD'(x"0974090a"),
RAM_WORD'(x"8106ff05"),
RAM_WORD'(x"06075351"),
RAM_WORD'(x"04000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"71715351"),
RAM_WORD'(x"04067383"),
RAM_WORD'(x"06098105"),
RAM_WORD'(x"8205832b"),
RAM_WORD'(x"0b2b0772"),
RAM_WORD'(x"fc060c51"),
RAM_WORD'(x"51040000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"72098105"),
RAM_WORD'(x"72050970"),
RAM_WORD'(x"81050906"),
RAM_WORD'(x"0a810653"),
RAM_WORD'(x"51040000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"72098105"),
RAM_WORD'(x"72050970"),
RAM_WORD'(x"81050906"),
RAM_WORD'(x"0a098106"),
RAM_WORD'(x"53510400"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"71098105"),
RAM_WORD'(x"52040000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"72720981"),
RAM_WORD'(x"05055351"),
RAM_WORD'(x"04000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"72097206"),
RAM_WORD'(x"73730906"),
RAM_WORD'(x"07535104"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"71fc0608"),
RAM_WORD'(x"72830609"),
RAM_WORD'(x"81058305"),
RAM_WORD'(x"1010102a"),
RAM_WORD'(x"81ff0652"),
RAM_WORD'(x"04000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"71fc0608"),
RAM_WORD'(x"0b0b8180"),
RAM_WORD'(x"80738306"),
RAM_WORD'(x"10100508"),
RAM_WORD'(x"060b0b0b"),
RAM_WORD'(x"88a90400"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"0b0b0b89"),
RAM_WORD'(x"85040000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"0b0b0b88"),
RAM_WORD'(x"df040000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"72097081"),
RAM_WORD'(x"0509060a"),
RAM_WORD'(x"8106ff05"),
RAM_WORD'(x"70547106"),
RAM_WORD'(x"73097274"),
RAM_WORD'(x"05ff0506"),
RAM_WORD'(x"07515151"),
RAM_WORD'(x"04000000"),
RAM_WORD'(x"72097081"),
RAM_WORD'(x"0509060a"),
RAM_WORD'(x"098106ff"),
RAM_WORD'(x"05705471"),
RAM_WORD'(x"06730972"),
RAM_WORD'(x"7405ff05"),
RAM_WORD'(x"06075151"),
RAM_WORD'(x"51040000"),
RAM_WORD'(x"05ff0504"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"810b0b0b"),
RAM_WORD'(x"8180900c"),
RAM_WORD'(x"51040000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"71810552"),
RAM_WORD'(x"04000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"02840572"),
RAM_WORD'(x"05520400"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"717105ff"),
RAM_WORD'(x"05715351"),
RAM_WORD'(x"04000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"81fb3fae"),
RAM_WORD'(x"9e3f0410"),
RAM_WORD'(x"10101010"),
RAM_WORD'(x"10101010"),
RAM_WORD'(x"10101010"),
RAM_WORD'(x"10101010"),
RAM_WORD'(x"10101010"),
RAM_WORD'(x"10101010"),
RAM_WORD'(x"10101010"),
RAM_WORD'(x"10105351"),
RAM_WORD'(x"047381ff"),
RAM_WORD'(x"06738306"),
RAM_WORD'(x"09810583"),
RAM_WORD'(x"05101010"),
RAM_WORD'(x"2b0772fc"),
RAM_WORD'(x"060c5151"),
RAM_WORD'(x"043c0472"),
RAM_WORD'(x"72807281"),
RAM_WORD'(x"06ff0509"),
RAM_WORD'(x"72060571"),
RAM_WORD'(x"1052720a"),
RAM_WORD'(x"100a5372"),
RAM_WORD'(x"ed385151"),
RAM_WORD'(x"53510481"),
RAM_WORD'(x"90980881"),
RAM_WORD'(x"909c0881"),
RAM_WORD'(x"90a00875"),
RAM_WORD'(x"759c912d"),
RAM_WORD'(x"50508190"),
RAM_WORD'(x"98085681"),
RAM_WORD'(x"90a00c81"),
RAM_WORD'(x"909c0c81"),
RAM_WORD'(x"90980c51"),
RAM_WORD'(x"04819098"),
RAM_WORD'(x"0881909c"),
RAM_WORD'(x"088190a0"),
RAM_WORD'(x"0875759a"),
RAM_WORD'(x"a52d5050"),
RAM_WORD'(x"81909808"),
RAM_WORD'(x"568190a0"),
RAM_WORD'(x"0c81909c"),
RAM_WORD'(x"0c819098"),
RAM_WORD'(x"0c510481"),
RAM_WORD'(x"90980881"),
RAM_WORD'(x"909c0881"),
RAM_WORD'(x"90a008b6"),
RAM_WORD'(x"a02d8190"),
RAM_WORD'(x"a00c8190"),
RAM_WORD'(x"9c0c8190"),
RAM_WORD'(x"980c04fc"),
RAM_WORD'(x"3d0d818f"),
RAM_WORD'(x"fc335170"),
RAM_WORD'(x"a7388180"),
RAM_WORD'(x"9c087008"),
RAM_WORD'(x"52527080"),
RAM_WORD'(x"2e943884"),
RAM_WORD'(x"1281809c"),
RAM_WORD'(x"0c702d81"),
RAM_WORD'(x"809c0870"),
RAM_WORD'(x"08525270"),
RAM_WORD'(x"ee38810b"),
RAM_WORD'(x"818ffc34"),
RAM_WORD'(x"8c3d0d04"),
RAM_WORD'(x"04803d0d"),
RAM_WORD'(x"0b0b818f"),
RAM_WORD'(x"f408802e"),
RAM_WORD'(x"8e380b0b"),
RAM_WORD'(x"0b0b800b"),
RAM_WORD'(x"802e0981"),
RAM_WORD'(x"06853888"),
RAM_WORD'(x"3d0d040b"),
RAM_WORD'(x"0b818ff4"),
RAM_WORD'(x"510b0b0b"),
RAM_WORD'(x"f5da3f88"),
RAM_WORD'(x"3d0d0404"),
RAM_WORD'(x"f83d0d02"),
RAM_WORD'(x"93053353"),
RAM_WORD'(x"728a2e9d"),
RAM_WORD'(x"38819080"),
RAM_WORD'(x"08527108"),
RAM_WORD'(x"70882a81"),
RAM_WORD'(x"32708106"),
RAM_WORD'(x"51515170"),
RAM_WORD'(x"f1387272"),
RAM_WORD'(x"0c903d0d"),
RAM_WORD'(x"04819080"),
RAM_WORD'(x"08527108"),
RAM_WORD'(x"70882a81"),
RAM_WORD'(x"32708106"),
RAM_WORD'(x"51515170"),
RAM_WORD'(x"f1388d72"),
RAM_WORD'(x"0c710870"),
RAM_WORD'(x"882a8132"),
RAM_WORD'(x"70810651"),
RAM_WORD'(x"515170c2"),
RAM_WORD'(x"38d039fe"),
RAM_WORD'(x"e03d0d81"),
RAM_WORD'(x"ac3d7070"),
RAM_WORD'(x"84055208"),
RAM_WORD'(x"8aac5c55"),
RAM_WORD'(x"818c3d5e"),
RAM_WORD'(x"5c807470"),
RAM_WORD'(x"81055633"),
RAM_WORD'(x"755b5458"),
RAM_WORD'(x"72782e80"),
RAM_WORD'(x"c138b83d"),
RAM_WORD'(x"5b72a52e"),
RAM_WORD'(x"09810680"),
RAM_WORD'(x"c8387870"),
RAM_WORD'(x"81055a33"),
RAM_WORD'(x"537280e4"),
RAM_WORD'(x"2e81b938"),
RAM_WORD'(x"7280e424"),
RAM_WORD'(x"80c93872"),
RAM_WORD'(x"80e32ea4"),
RAM_WORD'(x"388052a5"),
RAM_WORD'(x"51792d80"),
RAM_WORD'(x"52725179"),
RAM_WORD'(x"2d821858"),
RAM_WORD'(x"78708105"),
RAM_WORD'(x"5a335372"),
RAM_WORD'(x"c4387781"),
RAM_WORD'(x"90980c81"),
RAM_WORD'(x"a83d0d04"),
RAM_WORD'(x"7b841d83"),
RAM_WORD'(x"1233555d"),
RAM_WORD'(x"56805272"),
RAM_WORD'(x"51792d81"),
RAM_WORD'(x"18797081"),
RAM_WORD'(x"055b3354"),
RAM_WORD'(x"5872ff9d"),
RAM_WORD'(x"38d83972"),
RAM_WORD'(x"80f32e09"),
RAM_WORD'(x"8106ffb5"),
RAM_WORD'(x"387b841d"),
RAM_WORD'(x"7108585d"),
RAM_WORD'(x"54807633"),
RAM_WORD'(x"58557675"),
RAM_WORD'(x"2e8d3881"),
RAM_WORD'(x"15701770"),
RAM_WORD'(x"33555855"),
RAM_WORD'(x"72f538ff"),
RAM_WORD'(x"15548075"),
RAM_WORD'(x"25ff9d38"),
RAM_WORD'(x"75708105"),
RAM_WORD'(x"57335380"),
RAM_WORD'(x"52725179"),
RAM_WORD'(x"2d811874"),
RAM_WORD'(x"ff165656"),
RAM_WORD'(x"58807525"),
RAM_WORD'(x"ff823875"),
RAM_WORD'(x"70810557"),
RAM_WORD'(x"33538052"),
RAM_WORD'(x"7251792d"),
RAM_WORD'(x"811874ff"),
RAM_WORD'(x"16565658"),
RAM_WORD'(x"748024cc"),
RAM_WORD'(x"38fee539"),
RAM_WORD'(x"7b841d71"),
RAM_WORD'(x"08555d55"),
RAM_WORD'(x"80732480"),
RAM_WORD'(x"f838727d"),
RAM_WORD'(x"7c565855"),
RAM_WORD'(x"80567276"),
RAM_WORD'(x"2e098106"),
RAM_WORD'(x"b638b07b"),
RAM_WORD'(x"3402b505"),
RAM_WORD'(x"547a742e"),
RAM_WORD'(x"9738ff14"),
RAM_WORD'(x"54733377"),
RAM_WORD'(x"70810559"),
RAM_WORD'(x"34811656"),
RAM_WORD'(x"7a742e09"),
RAM_WORD'(x"8106eb38"),
RAM_WORD'(x"80773475"),
RAM_WORD'(x"7dff1256"),
RAM_WORD'(x"57557480"),
RAM_WORD'(x"24fef938"),
RAM_WORD'(x"fe92398a"),
RAM_WORD'(x"7536b6e4"),
RAM_WORD'(x"05537233"),
RAM_WORD'(x"74708105"),
RAM_WORD'(x"56348a75"),
RAM_WORD'(x"35557480"),
RAM_WORD'(x"2effba38"),
RAM_WORD'(x"8a7536b6"),
RAM_WORD'(x"e4055372"),
RAM_WORD'(x"33747081"),
RAM_WORD'(x"0556348a"),
RAM_WORD'(x"75355574"),
RAM_WORD'(x"d238ffa1"),
RAM_WORD'(x"39723053"),
RAM_WORD'(x"ff8439fe"),
RAM_WORD'(x"f83d0db0"),
RAM_WORD'(x"5192df3f"),
RAM_WORD'(x"81909808"),
RAM_WORD'(x"81debc0c"),
RAM_WORD'(x"b05192d2"),
RAM_WORD'(x"3f819098"),
RAM_WORD'(x"0881decc"),
RAM_WORD'(x"0c81debc"),
RAM_WORD'(x"08819098"),
RAM_WORD'(x"080c800b"),
RAM_WORD'(x"81909808"),
RAM_WORD'(x"84050c82"),
RAM_WORD'(x"0b819098"),
RAM_WORD'(x"0888050c"),
RAM_WORD'(x"a80b8190"),
RAM_WORD'(x"98088c05"),
RAM_WORD'(x"0c9f53b6"),
RAM_WORD'(x"f0528190"),
RAM_WORD'(x"98089005"),
RAM_WORD'(x"519ec03f"),
RAM_WORD'(x"80f03d5b"),
RAM_WORD'(x"9f53b790"),
RAM_WORD'(x"527a519e"),
RAM_WORD'(x"b23f8a0b"),
RAM_WORD'(x"819d840c"),
RAM_WORD'(x"bbdc51fc"),
RAM_WORD'(x"923fb7b0"),
RAM_WORD'(x"51fc8c3f"),
RAM_WORD'(x"bbdc51fc"),
RAM_WORD'(x"863fb252"),
RAM_WORD'(x"b7e051fb"),
RAM_WORD'(x"fe3f8180"),
RAM_WORD'(x"a0085581"),
RAM_WORD'(x"750c8275"),
RAM_WORD'(x"0c740881"),
RAM_WORD'(x"90940c81"),
RAM_WORD'(x"0b80d43d"),
RAM_WORD'(x"80d03d42"),
RAM_WORD'(x"405a80c1"),
RAM_WORD'(x"0b81dec4"),
RAM_WORD'(x"34810b81"),
RAM_WORD'(x"e09c0c80"),
RAM_WORD'(x"c20b81de"),
RAM_WORD'(x"c8348242"),
RAM_WORD'(x"835e9f53"),
RAM_WORD'(x"b890527e"),
RAM_WORD'(x"519dd43f"),
RAM_WORD'(x"81438058"),
RAM_WORD'(x"820b81de"),
RAM_WORD'(x"c4330288"),
RAM_WORD'(x"0580cf05"),
RAM_WORD'(x"58585574"),
RAM_WORD'(x"1b703377"),
RAM_WORD'(x"33435154"),
RAM_WORD'(x"73612e87"),
RAM_WORD'(x"fe3880c1"),
RAM_WORD'(x"0b811681"),
RAM_WORD'(x"1858565c"),
RAM_WORD'(x"827525e3"),
RAM_WORD'(x"387681de"),
RAM_WORD'(x"c4347b80"),
RAM_WORD'(x"d22e9238"),
RAM_WORD'(x"7e527a51"),
RAM_WORD'(x"9eea3f80"),
RAM_WORD'(x"0b819098"),
RAM_WORD'(x"082587ce"),
RAM_WORD'(x"387781e0"),
RAM_WORD'(x"9c0c6170"),
RAM_WORD'(x"56567583"),
RAM_WORD'(x"25953881"),
RAM_WORD'(x"16548515"),
RAM_WORD'(x"74758117"),
RAM_WORD'(x"57575759"),
RAM_WORD'(x"837624f2"),
RAM_WORD'(x"38754285"),
RAM_WORD'(x"1670822b"),
RAM_WORD'(x"81ded411"),
RAM_WORD'(x"707c7170"),
RAM_WORD'(x"8405530c"),
RAM_WORD'(x"7c710c44"),
RAM_WORD'(x"7280f812"),
RAM_WORD'(x"0c577186"),
RAM_WORD'(x"19595759"),
RAM_WORD'(x"57767624"),
RAM_WORD'(x"9b3876b3"),
RAM_WORD'(x"29822b81"),
RAM_WORD'(x"90a81151"),
RAM_WORD'(x"54767470"),
RAM_WORD'(x"8405560c"),
RAM_WORD'(x"81155575"),
RAM_WORD'(x"7525f238"),
RAM_WORD'(x"7681cc29"),
RAM_WORD'(x"8190a805"),
RAM_WORD'(x"fc110881"),
RAM_WORD'(x"05fc120c"),
RAM_WORD'(x"81ded419"),
RAM_WORD'(x"089fa012"),
RAM_WORD'(x"0c56850b"),
RAM_WORD'(x"81dec00c"),
RAM_WORD'(x"81decc08"),
RAM_WORD'(x"70085755"),
RAM_WORD'(x"b0537452"),
RAM_WORD'(x"75519bf3"),
RAM_WORD'(x"3f850b8c"),
RAM_WORD'(x"160c850b"),
RAM_WORD'(x"8c170c74"),
RAM_WORD'(x"08760c81"),
RAM_WORD'(x"decc0854"),
RAM_WORD'(x"73802e8a"),
RAM_WORD'(x"38730876"),
RAM_WORD'(x"0c81decc"),
RAM_WORD'(x"085481de"),
RAM_WORD'(x"c0088c05"),
RAM_WORD'(x"8c150c84"),
RAM_WORD'(x"16085776"),
RAM_WORD'(x"86c23886"),
RAM_WORD'(x"0b8c170c"),
RAM_WORD'(x"88150888"),
RAM_WORD'(x"17565473"),
RAM_WORD'(x"822e86c8"),
RAM_WORD'(x"38835873"),
RAM_WORD'(x"812e86d7"),
RAM_WORD'(x"38817426"),
RAM_WORD'(x"86dc3873"),
RAM_WORD'(x"822e86b4"),
RAM_WORD'(x"3873842e"),
RAM_WORD'(x"85ff3877"),
RAM_WORD'(x"750c81de"),
RAM_WORD'(x"cc087008"),
RAM_WORD'(x"770c578c"),
RAM_WORD'(x"16088c05"),
RAM_WORD'(x"8c170c80"),
RAM_WORD'(x"c10b81de"),
RAM_WORD'(x"c8335656"),
RAM_WORD'(x"7481ff06"),
RAM_WORD'(x"41756126"),
RAM_WORD'(x"a2388054"),
RAM_WORD'(x"7580c32e"),
RAM_WORD'(x"85bc3873"),
RAM_WORD'(x"632e86b1"),
RAM_WORD'(x"38811670"),
RAM_WORD'(x"81ff0657"),
RAM_WORD'(x"547481ff"),
RAM_WORD'(x"06416076"),
RAM_WORD'(x"27e0387d"),
RAM_WORD'(x"62297971"),
RAM_WORD'(x"35704471"),
RAM_WORD'(x"7b317087"),
RAM_WORD'(x"2972315b"),
RAM_WORD'(x"578a0581"),
RAM_WORD'(x"dec43381"),
RAM_WORD'(x"dec0085a"),
RAM_WORD'(x"52555675"),
RAM_WORD'(x"80c12e86"),
RAM_WORD'(x"9c387cf7"),
RAM_WORD'(x"38811a5a"),
RAM_WORD'(x"b27a25fc"),
RAM_WORD'(x"a5388180"),
RAM_WORD'(x"a0085c82"),
RAM_WORD'(x"7c0c7b08"),
RAM_WORD'(x"7081deb8"),
RAM_WORD'(x"0c52b8b0"),
RAM_WORD'(x"51f7f03f"),
RAM_WORD'(x"81909408"),
RAM_WORD'(x"52b8c051"),
RAM_WORD'(x"f7e53fb8"),
RAM_WORD'(x"d051f7df"),
RAM_WORD'(x"3fbbdc51"),
RAM_WORD'(x"f7d93f81"),
RAM_WORD'(x"deb80881"),
RAM_WORD'(x"90940831"),
RAM_WORD'(x"70819090"),
RAM_WORD'(x"0cb27135"),
RAM_WORD'(x"8190880c"),
RAM_WORD'(x"70bd84c0"),
RAM_WORD'(x"3570b229"),
RAM_WORD'(x"81908c0c"),
RAM_WORD'(x"8ddd7183"),
RAM_WORD'(x"86d02935"),
RAM_WORD'(x"81ded00c"),
RAM_WORD'(x"57b8e052"),
RAM_WORD'(x"5df7a43f"),
RAM_WORD'(x"81908808"),
RAM_WORD'(x"52b8cc51"),
RAM_WORD'(x"f7993fb8"),
RAM_WORD'(x"f051f793"),
RAM_WORD'(x"3f81908c"),
RAM_WORD'(x"0852b980"),
RAM_WORD'(x"51f7883f"),
RAM_WORD'(x"81ded008"),
RAM_WORD'(x"52b98851"),
RAM_WORD'(x"f6fd3fbb"),
RAM_WORD'(x"dc51f6f7"),
RAM_WORD'(x"3fb99c51"),
RAM_WORD'(x"f6f13fbb"),
RAM_WORD'(x"dc51f6eb"),
RAM_WORD'(x"3f81dec0"),
RAM_WORD'(x"0852b9d4"),
RAM_WORD'(x"51f6e03f"),
RAM_WORD'(x"8552b9f0"),
RAM_WORD'(x"51f6d83f"),
RAM_WORD'(x"81e09c08"),
RAM_WORD'(x"52ba8c51"),
RAM_WORD'(x"f6cd3f81"),
RAM_WORD'(x"52b9f051"),
RAM_WORD'(x"f6c53f81"),
RAM_WORD'(x"dec43352"),
RAM_WORD'(x"baa851f6"),
RAM_WORD'(x"ba3f80c1"),
RAM_WORD'(x"52bac451"),
RAM_WORD'(x"f6b13f81"),
RAM_WORD'(x"dec83352"),
RAM_WORD'(x"bae051f6"),
RAM_WORD'(x"a63f80c2"),
RAM_WORD'(x"52bac451"),
RAM_WORD'(x"f69d3f81"),
RAM_WORD'(x"def40852"),
RAM_WORD'(x"bafc51f6"),
RAM_WORD'(x"923f8752"),
RAM_WORD'(x"b9f051f6"),
RAM_WORD'(x"8a3f819d"),
RAM_WORD'(x"840852bb"),
RAM_WORD'(x"9851f5ff"),
RAM_WORD'(x"3fbbb451"),
RAM_WORD'(x"f5f93fbb"),
RAM_WORD'(x"e051f5f3"),
RAM_WORD'(x"3f81decc"),
RAM_WORD'(x"08700853"),
RAM_WORD'(x"55bbec51"),
RAM_WORD'(x"f5e53fbc"),
RAM_WORD'(x"8851f5df"),
RAM_WORD'(x"3f81decc"),
RAM_WORD'(x"08841108"),
RAM_WORD'(x"535ebcbc"),
RAM_WORD'(x"51f5d03f"),
RAM_WORD'(x"8052b9f0"),
RAM_WORD'(x"51f5c83f"),
RAM_WORD'(x"81decc08"),
RAM_WORD'(x"88110853"),
RAM_WORD'(x"54bcd851"),
RAM_WORD'(x"f5b93f82"),
RAM_WORD'(x"52b9f051"),
RAM_WORD'(x"f5b13f81"),
RAM_WORD'(x"decc088c"),
RAM_WORD'(x"11085341"),
RAM_WORD'(x"bcf451f5"),
RAM_WORD'(x"a23f9152"),
RAM_WORD'(x"b9f051f5"),
RAM_WORD'(x"9a3f81de"),
RAM_WORD'(x"cc089005"),
RAM_WORD'(x"52bd9051"),
RAM_WORD'(x"f58d3fbd"),
RAM_WORD'(x"ac51f587"),
RAM_WORD'(x"3fbde451"),
RAM_WORD'(x"f5813f81"),
RAM_WORD'(x"debc0870"),
RAM_WORD'(x"085357bb"),
RAM_WORD'(x"ec51f4f3"),
RAM_WORD'(x"3fbdf851"),
RAM_WORD'(x"f4ed3f81"),
RAM_WORD'(x"debc0884"),
RAM_WORD'(x"11085340"),
RAM_WORD'(x"bcbc51f4"),
RAM_WORD'(x"de3f8052"),
RAM_WORD'(x"b9f051f4"),
RAM_WORD'(x"d63f81de"),
RAM_WORD'(x"bc088811"),
RAM_WORD'(x"08535cbc"),
RAM_WORD'(x"d851f4c7"),
RAM_WORD'(x"3f8152b9"),
RAM_WORD'(x"f051f4bf"),
RAM_WORD'(x"3f81debc"),
RAM_WORD'(x"088c1108"),
RAM_WORD'(x"535abcf4"),
RAM_WORD'(x"51f4b03f"),
RAM_WORD'(x"9252b9f0"),
RAM_WORD'(x"51f4a83f"),
RAM_WORD'(x"81debc08"),
RAM_WORD'(x"900552bd"),
RAM_WORD'(x"9051f49b"),
RAM_WORD'(x"3fbdac51"),
RAM_WORD'(x"f4953f61"),
RAM_WORD'(x"52beb851"),
RAM_WORD'(x"f48d3f85"),
RAM_WORD'(x"52b9f051"),
RAM_WORD'(x"f4853f77"),
RAM_WORD'(x"52bed451"),
RAM_WORD'(x"f3fd3f8d"),
RAM_WORD'(x"52b9f051"),
RAM_WORD'(x"f3f53f78"),
RAM_WORD'(x"52bef051"),
RAM_WORD'(x"f3ed3f87"),
RAM_WORD'(x"52b9f051"),
RAM_WORD'(x"f3e53f62"),
RAM_WORD'(x"52bf8c51"),
RAM_WORD'(x"f3dd3f81"),
RAM_WORD'(x"52b9f051"),
RAM_WORD'(x"f3d53f7a"),
RAM_WORD'(x"52bfa851"),
RAM_WORD'(x"f3cd3fbf"),
RAM_WORD'(x"c451f3c7"),
RAM_WORD'(x"3f7e520b"),
RAM_WORD'(x"bffc51f3"),
RAM_WORD'(x"be3f80c0"),
RAM_WORD'(x"9851f3b7"),
RAM_WORD'(x"3fbbdc51"),
RAM_WORD'(x"f3b13f80"),
RAM_WORD'(x"0b819098"),
RAM_WORD'(x"0c81903d"),
RAM_WORD'(x"0d048158"),
RAM_WORD'(x"f8af3973"),
RAM_WORD'(x"57827525"),
RAM_WORD'(x"f7ed38f8"),
RAM_WORD'(x"88397581"),
RAM_WORD'(x"dec43481"),
RAM_WORD'(x"5473632e"),
RAM_WORD'(x"098106fa"),
RAM_WORD'(x"bc3880e9"),
RAM_WORD'(x"3982750c"),
RAM_WORD'(x"81decc08"),
RAM_WORD'(x"7008770c"),
RAM_WORD'(x"578c1608"),
RAM_WORD'(x"8c058c17"),
RAM_WORD'(x"0cfa8039"),
RAM_WORD'(x"740858b0"),
RAM_WORD'(x"53775274"),
RAM_WORD'(x"5194f43f"),
RAM_WORD'(x"80c10b81"),
RAM_WORD'(x"dec83356"),
RAM_WORD'(x"56f9f139"),
RAM_WORD'(x"81750c81"),
RAM_WORD'(x"decc0870"),
RAM_WORD'(x"08770c57"),
RAM_WORD'(x"8c16088c"),
RAM_WORD'(x"058c170c"),
RAM_WORD'(x"f9d13980"),
RAM_WORD'(x"e40b81de"),
RAM_WORD'(x"c00825f9"),
RAM_WORD'(x"b2387675"),
RAM_WORD'(x"0c81decc"),
RAM_WORD'(x"08700877"),
RAM_WORD'(x"0c578c16"),
RAM_WORD'(x"088c058c"),
RAM_WORD'(x"170cf9af"),
RAM_WORD'(x"3980439f"),
RAM_WORD'(x"5380c0d0"),
RAM_WORD'(x"527e5194"),
RAM_WORD'(x"a23f797a"),
RAM_WORD'(x"81dec00c"),
RAM_WORD'(x"81dec833"),
RAM_WORD'(x"81187081"),
RAM_WORD'(x"ff065956"),
RAM_WORD'(x"565ef9b5"),
RAM_WORD'(x"39ff1470"),
RAM_WORD'(x"7831610c"),
RAM_WORD'(x"5d800b81"),
RAM_WORD'(x"1b5b5db2"),
RAM_WORD'(x"7a25f682"),
RAM_WORD'(x"38f9db39"),
RAM_WORD'(x"f43d0d80"),
RAM_WORD'(x"c0f40b81"),
RAM_WORD'(x"80805454"),
RAM_WORD'(x"73708405"),
RAM_WORD'(x"55087370"),
RAM_WORD'(x"8405550c"),
RAM_WORD'(x"818ff473"),
RAM_WORD'(x"26ee3880"),
RAM_WORD'(x"d0f80b81"),
RAM_WORD'(x"8ff45454"),
RAM_WORD'(x"72818ff8"),
RAM_WORD'(x"27943873"),
RAM_WORD'(x"70840555"),
RAM_WORD'(x"08737084"),
RAM_WORD'(x"05550c81"),
RAM_WORD'(x"8ff87326"),
RAM_WORD'(x"ee388280"),
RAM_WORD'(x"800b8190"),
RAM_WORD'(x"800c8380"),
RAM_WORD'(x"800b8190"),
RAM_WORD'(x"840c0b0b"),
RAM_WORD'(x"0bb6d40b"),
RAM_WORD'(x"818ff80c"),
RAM_WORD'(x"ee823f81"),
RAM_WORD'(x"80ac5281"),
RAM_WORD'(x"51f3fc3f"),
RAM_WORD'(x"81909808"),
RAM_WORD'(x"5185b73f"),
RAM_WORD'(x"803d0d81"),
RAM_WORD'(x"80a80813"),
RAM_WORD'(x"708180a8"),
RAM_WORD'(x"0c819098"),
RAM_WORD'(x"0c883d0d"),
RAM_WORD'(x"048190a4"),
RAM_WORD'(x"08028190"),
RAM_WORD'(x"a40ce43d"),
RAM_WORD'(x"0d800b81"),
RAM_WORD'(x"90a408fc"),
RAM_WORD'(x"050c8190"),
RAM_WORD'(x"a4088805"),
RAM_WORD'(x"088025b9"),
RAM_WORD'(x"388190a4"),
RAM_WORD'(x"08880508"),
RAM_WORD'(x"308190a4"),
RAM_WORD'(x"0888050c"),
RAM_WORD'(x"800b8190"),
RAM_WORD'(x"a408f405"),
RAM_WORD'(x"0c8190a4"),
RAM_WORD'(x"08fc0508"),
RAM_WORD'(x"8a38810b"),
RAM_WORD'(x"8190a408"),
RAM_WORD'(x"f4050c81"),
RAM_WORD'(x"90a408f4"),
RAM_WORD'(x"05088190"),
RAM_WORD'(x"a408fc05"),
RAM_WORD'(x"0c8190a4"),
RAM_WORD'(x"088c0508"),
RAM_WORD'(x"8025b938"),
RAM_WORD'(x"8190a408"),
RAM_WORD'(x"8c050830"),
RAM_WORD'(x"8190a408"),
RAM_WORD'(x"8c050c80"),
RAM_WORD'(x"0b8190a4"),
RAM_WORD'(x"08f0050c"),
RAM_WORD'(x"8190a408"),
RAM_WORD'(x"fc05088a"),
RAM_WORD'(x"38810b81"),
RAM_WORD'(x"90a408f0"),
RAM_WORD'(x"050c8190"),
RAM_WORD'(x"a408f005"),
RAM_WORD'(x"088190a4"),
RAM_WORD'(x"08fc050c"),
RAM_WORD'(x"80538190"),
RAM_WORD'(x"a4088c05"),
RAM_WORD'(x"08528190"),
RAM_WORD'(x"a4088805"),
RAM_WORD'(x"085181df"),
RAM_WORD'(x"3f819098"),
RAM_WORD'(x"08708190"),
RAM_WORD'(x"a408f805"),
RAM_WORD'(x"0c548190"),
RAM_WORD'(x"a408fc05"),
RAM_WORD'(x"08802e90"),
RAM_WORD'(x"388190a4"),
RAM_WORD'(x"08f80508"),
RAM_WORD'(x"308190a4"),
RAM_WORD'(x"08f8050c"),
RAM_WORD'(x"8190a408"),
RAM_WORD'(x"f8050870"),
RAM_WORD'(x"8190980c"),
RAM_WORD'(x"54a43d0d"),
RAM_WORD'(x"8190a40c"),
RAM_WORD'(x"048190a4"),
RAM_WORD'(x"08028190"),
RAM_WORD'(x"a40cec3d"),
RAM_WORD'(x"0d800b81"),
RAM_WORD'(x"90a408fc"),
RAM_WORD'(x"050c8190"),
RAM_WORD'(x"a4088805"),
RAM_WORD'(x"08802599"),
RAM_WORD'(x"388190a4"),
RAM_WORD'(x"08880508"),
RAM_WORD'(x"308190a4"),
RAM_WORD'(x"0888050c"),
RAM_WORD'(x"810b8190"),
RAM_WORD'(x"a408fc05"),
RAM_WORD'(x"0c8190a4"),
RAM_WORD'(x"088c0508"),
RAM_WORD'(x"80259038"),
RAM_WORD'(x"8190a408"),
RAM_WORD'(x"8c050830"),
RAM_WORD'(x"8190a408"),
RAM_WORD'(x"8c050c81"),
RAM_WORD'(x"538190a4"),
RAM_WORD'(x"088c0508"),
RAM_WORD'(x"528190a4"),
RAM_WORD'(x"08880508"),
RAM_WORD'(x"51bd3f81"),
RAM_WORD'(x"90980870"),
RAM_WORD'(x"8190a408"),
RAM_WORD'(x"f8050c54"),
RAM_WORD'(x"8190a408"),
RAM_WORD'(x"fc050880"),
RAM_WORD'(x"2e903881"),
RAM_WORD'(x"90a408f8"),
RAM_WORD'(x"05083081"),
RAM_WORD'(x"90a408f8"),
RAM_WORD'(x"050c8190"),
RAM_WORD'(x"a408f805"),
RAM_WORD'(x"08708190"),
RAM_WORD'(x"980c549c"),
RAM_WORD'(x"3d0d8190"),
RAM_WORD'(x"a40c0481"),
RAM_WORD'(x"90a40802"),
RAM_WORD'(x"8190a40c"),
RAM_WORD'(x"f43d0d81"),
RAM_WORD'(x"0b8190a4"),
RAM_WORD'(x"08fc050c"),
RAM_WORD'(x"800b8190"),
RAM_WORD'(x"a408f805"),
RAM_WORD'(x"0c8190a4"),
RAM_WORD'(x"088c0508"),
RAM_WORD'(x"8190a408"),
RAM_WORD'(x"88050827"),
RAM_WORD'(x"b9388190"),
RAM_WORD'(x"a408fc05"),
RAM_WORD'(x"08802eae"),
RAM_WORD'(x"38800b81"),
RAM_WORD'(x"90a4088c"),
RAM_WORD'(x"050824a2"),
RAM_WORD'(x"388190a4"),
RAM_WORD'(x"088c0508"),
RAM_WORD'(x"108190a4"),
RAM_WORD'(x"088c050c"),
RAM_WORD'(x"8190a408"),
RAM_WORD'(x"fc050810"),
RAM_WORD'(x"8190a408"),
RAM_WORD'(x"fc050cff"),
RAM_WORD'(x"b8398190"),
RAM_WORD'(x"a408fc05"),
RAM_WORD'(x"08802e80"),
RAM_WORD'(x"e1388190"),
RAM_WORD'(x"a4088c05"),
RAM_WORD'(x"088190a4"),
RAM_WORD'(x"08880508"),
RAM_WORD'(x"26ad3881"),
RAM_WORD'(x"90a40888"),
RAM_WORD'(x"05088190"),
RAM_WORD'(x"a4088c05"),
RAM_WORD'(x"08318190"),
RAM_WORD'(x"a4088805"),
RAM_WORD'(x"0c8190a4"),
RAM_WORD'(x"08f80508"),
RAM_WORD'(x"8190a408"),
RAM_WORD'(x"fc050807"),
RAM_WORD'(x"8190a408"),
RAM_WORD'(x"f8050c81"),
RAM_WORD'(x"90a408fc"),
RAM_WORD'(x"0508812a"),
RAM_WORD'(x"8190a408"),
RAM_WORD'(x"fc050c81"),
RAM_WORD'(x"90a4088c"),
RAM_WORD'(x"0508812a"),
RAM_WORD'(x"8190a408"),
RAM_WORD'(x"8c050cff"),
RAM_WORD'(x"95398190"),
RAM_WORD'(x"a4089005"),
RAM_WORD'(x"08802e93"),
RAM_WORD'(x"388190a4"),
RAM_WORD'(x"08880508"),
RAM_WORD'(x"708190a4"),
RAM_WORD'(x"08f4050c"),
RAM_WORD'(x"51913981"),
RAM_WORD'(x"90a408f8"),
RAM_WORD'(x"05087081"),
RAM_WORD'(x"90a408f4"),
RAM_WORD'(x"050c5181"),
RAM_WORD'(x"90a408f4"),
RAM_WORD'(x"05088190"),
RAM_WORD'(x"980c943d"),
RAM_WORD'(x"0d8190a4"),
RAM_WORD'(x"0c04dc3d"),
RAM_WORD'(x"0d7b8180"),
RAM_WORD'(x"b00882c8"),
RAM_WORD'(x"11085a54"),
RAM_WORD'(x"5a77802e"),
RAM_WORD'(x"80da3881"),
RAM_WORD'(x"88188419"),
RAM_WORD'(x"08ff0581"),
RAM_WORD'(x"712b5955"),
RAM_WORD'(x"59807424"),
RAM_WORD'(x"80ea3880"),
RAM_WORD'(x"7424b538"),
RAM_WORD'(x"73822b78"),
RAM_WORD'(x"11880556"),
RAM_WORD'(x"56818019"),
RAM_WORD'(x"08770653"),
RAM_WORD'(x"72802eb6"),
RAM_WORD'(x"38781670"),
RAM_WORD'(x"08535379"),
RAM_WORD'(x"51740853"),
RAM_WORD'(x"722dff14"),
RAM_WORD'(x"fc17fc17"),
RAM_WORD'(x"79812c5a"),
RAM_WORD'(x"57575473"),
RAM_WORD'(x"8025d638"),
RAM_WORD'(x"77085877"),
RAM_WORD'(x"ffad3881"),
RAM_WORD'(x"80b00853"),
RAM_WORD'(x"bc1308a5"),
RAM_WORD'(x"38795195"),
RAM_WORD'(x"e03f7408"),
RAM_WORD'(x"53722dff"),
RAM_WORD'(x"14fc17fc"),
RAM_WORD'(x"1779812c"),
RAM_WORD'(x"5a575754"),
RAM_WORD'(x"738025ff"),
RAM_WORD'(x"a838d139"),
RAM_WORD'(x"8057ff93"),
RAM_WORD'(x"397251bc"),
RAM_WORD'(x"13085372"),
RAM_WORD'(x"2d795195"),
RAM_WORD'(x"b43ffc3d"),
RAM_WORD'(x"0d735281"),
RAM_WORD'(x"80b00851"),
RAM_WORD'(x"963f8c3d"),
RAM_WORD'(x"0d04fc3d"),
RAM_WORD'(x"0d735281"),
RAM_WORD'(x"80b00851"),
RAM_WORD'(x"90c13f8c"),
RAM_WORD'(x"3d0d04cc"),
RAM_WORD'(x"3d0d7f61"),
RAM_WORD'(x"8b1170f8"),
RAM_WORD'(x"065c5555"),
RAM_WORD'(x"5e729626"),
RAM_WORD'(x"83389059"),
RAM_WORD'(x"80792474"),
RAM_WORD'(x"7a260753"),
RAM_WORD'(x"80547274"),
RAM_WORD'(x"2e098106"),
RAM_WORD'(x"80cb387d"),
RAM_WORD'(x"518cf73f"),
RAM_WORD'(x"7883f726"),
RAM_WORD'(x"80c83878"),
RAM_WORD'(x"832a7010"),
RAM_WORD'(x"10108187"),
RAM_WORD'(x"ec058c11"),
RAM_WORD'(x"0859595a"),
RAM_WORD'(x"76782e83"),
RAM_WORD'(x"b2388417"),
RAM_WORD'(x"08fc0656"),
RAM_WORD'(x"8c170888"),
RAM_WORD'(x"1808718c"),
RAM_WORD'(x"120c8812"),
RAM_WORD'(x"0c587517"),
RAM_WORD'(x"84110881"),
RAM_WORD'(x"0784120c"),
RAM_WORD'(x"537d518c"),
RAM_WORD'(x"b63f8817"),
RAM_WORD'(x"54738190"),
RAM_WORD'(x"980cbc3d"),
RAM_WORD'(x"0d047889"),
RAM_WORD'(x"2a79832a"),
RAM_WORD'(x"5b537280"),
RAM_WORD'(x"2ebf3878"),
RAM_WORD'(x"862ab805"),
RAM_WORD'(x"5a847327"),
RAM_WORD'(x"b43880db"),
RAM_WORD'(x"135a9473"),
RAM_WORD'(x"27ab3878"),
RAM_WORD'(x"8c2a80ee"),
RAM_WORD'(x"055a80d4"),
RAM_WORD'(x"73279e38"),
RAM_WORD'(x"788f2a80"),
RAM_WORD'(x"f7055a82"),
RAM_WORD'(x"d4732791"),
RAM_WORD'(x"3878922a"),
RAM_WORD'(x"80fc055a"),
RAM_WORD'(x"8ad47327"),
RAM_WORD'(x"843880fe"),
RAM_WORD'(x"5a791010"),
RAM_WORD'(x"108187ec"),
RAM_WORD'(x"058c1108"),
RAM_WORD'(x"58557675"),
RAM_WORD'(x"2ea33884"),
RAM_WORD'(x"1708fc06"),
RAM_WORD'(x"707a3155"),
RAM_WORD'(x"56738f24"),
RAM_WORD'(x"88e53873"),
RAM_WORD'(x"8025fee4"),
RAM_WORD'(x"388c1708"),
RAM_WORD'(x"5776752e"),
RAM_WORD'(x"098106df"),
RAM_WORD'(x"38811a5a"),
RAM_WORD'(x"8187fc08"),
RAM_WORD'(x"57768187"),
RAM_WORD'(x"f42e82c0"),
RAM_WORD'(x"38841708"),
RAM_WORD'(x"fc06707a"),
RAM_WORD'(x"31555673"),
RAM_WORD'(x"8f2481f9"),
RAM_WORD'(x"388187f4"),
RAM_WORD'(x"0b818880"),
RAM_WORD'(x"0c8187f4"),
RAM_WORD'(x"0b8187fc"),
RAM_WORD'(x"0c738025"),
RAM_WORD'(x"feb03883"),
RAM_WORD'(x"ff762783"),
RAM_WORD'(x"e5387589"),
RAM_WORD'(x"2a76832a"),
RAM_WORD'(x"55537280"),
RAM_WORD'(x"2ebf3875"),
RAM_WORD'(x"862ab805"),
RAM_WORD'(x"54847327"),
RAM_WORD'(x"b43880db"),
RAM_WORD'(x"13549473"),
RAM_WORD'(x"27ab3875"),
RAM_WORD'(x"8c2a80ee"),
RAM_WORD'(x"055480d4"),
RAM_WORD'(x"73279e38"),
RAM_WORD'(x"758f2a80"),
RAM_WORD'(x"f7055482"),
RAM_WORD'(x"d4732791"),
RAM_WORD'(x"3875922a"),
RAM_WORD'(x"80fc0554"),
RAM_WORD'(x"8ad47327"),
RAM_WORD'(x"843880fe"),
RAM_WORD'(x"54731010"),
RAM_WORD'(x"108187ec"),
RAM_WORD'(x"05881108"),
RAM_WORD'(x"56587478"),
RAM_WORD'(x"2e86df38"),
RAM_WORD'(x"841508fc"),
RAM_WORD'(x"06537573"),
RAM_WORD'(x"278d3888"),
RAM_WORD'(x"15085574"),
RAM_WORD'(x"782e0981"),
RAM_WORD'(x"06ea388c"),
RAM_WORD'(x"15088187"),
RAM_WORD'(x"ec0b8405"),
RAM_WORD'(x"08718c1a"),
RAM_WORD'(x"0c76881a"),
RAM_WORD'(x"0c788813"),
RAM_WORD'(x"0c788c18"),
RAM_WORD'(x"0c5d5879"),
RAM_WORD'(x"53807a24"),
RAM_WORD'(x"83ec3872"),
RAM_WORD'(x"822c8171"),
RAM_WORD'(x"2b5c537a"),
RAM_WORD'(x"7c268198"),
RAM_WORD'(x"387b7b06"),
RAM_WORD'(x"537282f7"),
RAM_WORD'(x"3879fc06"),
RAM_WORD'(x"84055a7a"),
RAM_WORD'(x"10707d06"),
RAM_WORD'(x"545b7282"),
RAM_WORD'(x"e638841a"),
RAM_WORD'(x"5af13988"),
RAM_WORD'(x"178c1108"),
RAM_WORD'(x"58587678"),
RAM_WORD'(x"2e098106"),
RAM_WORD'(x"fcc03882"),
RAM_WORD'(x"1a5afdec"),
RAM_WORD'(x"39781779"),
RAM_WORD'(x"81078419"),
RAM_WORD'(x"0c708188"),
RAM_WORD'(x"800c7081"),
RAM_WORD'(x"87fc0c81"),
RAM_WORD'(x"87f40b8c"),
RAM_WORD'(x"120c8c11"),
RAM_WORD'(x"0888120c"),
RAM_WORD'(x"74810784"),
RAM_WORD'(x"120c7411"),
RAM_WORD'(x"75710c51"),
RAM_WORD'(x"537d5188"),
RAM_WORD'(x"e23f8817"),
RAM_WORD'(x"54fcaa39"),
RAM_WORD'(x"8187ec0b"),
RAM_WORD'(x"8405087a"),
RAM_WORD'(x"545c7980"),
RAM_WORD'(x"25fef838"),
RAM_WORD'(x"82e0397a"),
RAM_WORD'(x"097c0670"),
RAM_WORD'(x"8187ec0b"),
RAM_WORD'(x"84050c5c"),
RAM_WORD'(x"7a105b7a"),
RAM_WORD'(x"7c268538"),
RAM_WORD'(x"7a85c838"),
RAM_WORD'(x"8187ec0b"),
RAM_WORD'(x"88050870"),
RAM_WORD'(x"841208fc"),
RAM_WORD'(x"06707c31"),
RAM_WORD'(x"7c72268f"),
RAM_WORD'(x"72250757"),
RAM_WORD'(x"575c5d55"),
RAM_WORD'(x"72802e80"),
RAM_WORD'(x"e138797a"),
RAM_WORD'(x"168187e4"),
RAM_WORD'(x"081b9011"),
RAM_WORD'(x"5a55575b"),
RAM_WORD'(x"8187e008"),
RAM_WORD'(x"ff2e8838"),
RAM_WORD'(x"a08f13e0"),
RAM_WORD'(x"80065776"),
RAM_WORD'(x"527d5187"),
RAM_WORD'(x"eb3f8190"),
RAM_WORD'(x"98085481"),
RAM_WORD'(x"909808ff"),
RAM_WORD'(x"2e923881"),
RAM_WORD'(x"90980876"),
RAM_WORD'(x"27829938"),
RAM_WORD'(x"748187ec"),
RAM_WORD'(x"2e829138"),
RAM_WORD'(x"8187ec0b"),
RAM_WORD'(x"88050855"),
RAM_WORD'(x"841508fc"),
RAM_WORD'(x"06707a31"),
RAM_WORD'(x"7a72268f"),
RAM_WORD'(x"72250752"),
RAM_WORD'(x"55537283"),
RAM_WORD'(x"ee387479"),
RAM_WORD'(x"81078417"),
RAM_WORD'(x"0c791670"),
RAM_WORD'(x"8187ec0b"),
RAM_WORD'(x"88050c75"),
RAM_WORD'(x"81078412"),
RAM_WORD'(x"0c547e52"),
RAM_WORD'(x"5787903f"),
RAM_WORD'(x"881754fa"),
RAM_WORD'(x"d8397583"),
RAM_WORD'(x"2a705454"),
RAM_WORD'(x"80742481"),
RAM_WORD'(x"9b387282"),
RAM_WORD'(x"2c81712b"),
RAM_WORD'(x"8187f008"),
RAM_WORD'(x"07708187"),
RAM_WORD'(x"ec0b8405"),
RAM_WORD'(x"0c751010"),
RAM_WORD'(x"108187ec"),
RAM_WORD'(x"05881108"),
RAM_WORD'(x"585a5d53"),
RAM_WORD'(x"778c180c"),
RAM_WORD'(x"7488180c"),
RAM_WORD'(x"7688190c"),
RAM_WORD'(x"768c160c"),
RAM_WORD'(x"fced3979"),
RAM_WORD'(x"7a101010"),
RAM_WORD'(x"8187ec05"),
RAM_WORD'(x"7057595d"),
RAM_WORD'(x"8c150857"),
RAM_WORD'(x"76752ea3"),
RAM_WORD'(x"38841708"),
RAM_WORD'(x"fc06707a"),
RAM_WORD'(x"31555673"),
RAM_WORD'(x"8f2483d4"),
RAM_WORD'(x"38738025"),
RAM_WORD'(x"848b388c"),
RAM_WORD'(x"17085776"),
RAM_WORD'(x"752e0981"),
RAM_WORD'(x"06df3888"),
RAM_WORD'(x"15811b70"),
RAM_WORD'(x"8306555b"),
RAM_WORD'(x"5572c938"),
RAM_WORD'(x"7c830653"),
RAM_WORD'(x"72802efd"),
RAM_WORD'(x"b238ff1d"),
RAM_WORD'(x"f819595d"),
RAM_WORD'(x"88180878"),
RAM_WORD'(x"2eea38fd"),
RAM_WORD'(x"af39831a"),
RAM_WORD'(x"53fc9039"),
RAM_WORD'(x"83147082"),
RAM_WORD'(x"2c81712b"),
RAM_WORD'(x"8187f008"),
RAM_WORD'(x"07708187"),
RAM_WORD'(x"ec0b8405"),
RAM_WORD'(x"0c761010"),
RAM_WORD'(x"108187ec"),
RAM_WORD'(x"05881108"),
RAM_WORD'(x"595b5e51"),
RAM_WORD'(x"53fee139"),
RAM_WORD'(x"8187b008"),
RAM_WORD'(x"17588190"),
RAM_WORD'(x"9808762e"),
RAM_WORD'(x"81913881"),
RAM_WORD'(x"87e008ff"),
RAM_WORD'(x"2e83f438"),
RAM_WORD'(x"73763118"),
RAM_WORD'(x"8187b00c"),
RAM_WORD'(x"73870670"),
RAM_WORD'(x"57537280"),
RAM_WORD'(x"2e883888"),
RAM_WORD'(x"73317015"),
RAM_WORD'(x"55567614"),
RAM_WORD'(x"9fff06a0"),
RAM_WORD'(x"80713117"),
RAM_WORD'(x"70547f53"),
RAM_WORD'(x"575384f8"),
RAM_WORD'(x"3f819098"),
RAM_WORD'(x"08538190"),
RAM_WORD'(x"9808ff2e"),
RAM_WORD'(x"81a23881"),
RAM_WORD'(x"87b00816"),
RAM_WORD'(x"708187b0"),
RAM_WORD'(x"0c747581"),
RAM_WORD'(x"87ec0b88"),
RAM_WORD'(x"050c7476"),
RAM_WORD'(x"31187081"),
RAM_WORD'(x"07515556"),
RAM_WORD'(x"587b8187"),
RAM_WORD'(x"ec2e83a0"),
RAM_WORD'(x"38798f26"),
RAM_WORD'(x"82cf3881"),
RAM_WORD'(x"0b84150c"),
RAM_WORD'(x"841508fc"),
RAM_WORD'(x"06707a31"),
RAM_WORD'(x"7a72268f"),
RAM_WORD'(x"72250752"),
RAM_WORD'(x"55537280"),
RAM_WORD'(x"2efcf338"),
RAM_WORD'(x"80dd3981"),
RAM_WORD'(x"9098089f"),
RAM_WORD'(x"ff065372"),
RAM_WORD'(x"fee53877"),
RAM_WORD'(x"8187b00c"),
RAM_WORD'(x"8187ec0b"),
RAM_WORD'(x"8805087b"),
RAM_WORD'(x"18810784"),
RAM_WORD'(x"120c5581"),
RAM_WORD'(x"87dc0878"),
RAM_WORD'(x"27863877"),
RAM_WORD'(x"8187dc0c"),
RAM_WORD'(x"8187d808"),
RAM_WORD'(x"7827fca4"),
RAM_WORD'(x"38778187"),
RAM_WORD'(x"d80c8415"),
RAM_WORD'(x"08fc0670"),
RAM_WORD'(x"7a317a72"),
RAM_WORD'(x"268f7225"),
RAM_WORD'(x"07525553"),
RAM_WORD'(x"72802efc"),
RAM_WORD'(x"9d388839"),
RAM_WORD'(x"80745456"),
RAM_WORD'(x"fed9397d"),
RAM_WORD'(x"5183bc3f"),
RAM_WORD'(x"800b8190"),
RAM_WORD'(x"980cbc3d"),
RAM_WORD'(x"0d047353"),
RAM_WORD'(x"807424a9"),
RAM_WORD'(x"3872822c"),
RAM_WORD'(x"81712b81"),
RAM_WORD'(x"87f00807"),
RAM_WORD'(x"708187ec"),
RAM_WORD'(x"0b84050c"),
RAM_WORD'(x"5d53778c"),
RAM_WORD'(x"180c7488"),
RAM_WORD'(x"180c7688"),
RAM_WORD'(x"190c768c"),
RAM_WORD'(x"160cf9a7"),
RAM_WORD'(x"39831470"),
RAM_WORD'(x"822c8171"),
RAM_WORD'(x"2b8187f0"),
RAM_WORD'(x"08077081"),
RAM_WORD'(x"87ec0b84"),
RAM_WORD'(x"050c5e51"),
RAM_WORD'(x"53d4397b"),
RAM_WORD'(x"7b065372"),
RAM_WORD'(x"fc993884"),
RAM_WORD'(x"1a7b105c"),
RAM_WORD'(x"5af139ff"),
RAM_WORD'(x"1a811151"),
RAM_WORD'(x"5af7a939"),
RAM_WORD'(x"78177981"),
RAM_WORD'(x"0784190c"),
RAM_WORD'(x"8c180888"),
RAM_WORD'(x"1908718c"),
RAM_WORD'(x"120c8812"),
RAM_WORD'(x"0c597081"),
RAM_WORD'(x"88800c70"),
RAM_WORD'(x"8187fc0c"),
RAM_WORD'(x"8187f40b"),
RAM_WORD'(x"8c120c8c"),
RAM_WORD'(x"11088812"),
RAM_WORD'(x"0c748107"),
RAM_WORD'(x"84120c74"),
RAM_WORD'(x"1175710c"),
RAM_WORD'(x"5153f9ad"),
RAM_WORD'(x"39751784"),
RAM_WORD'(x"11088107"),
RAM_WORD'(x"84120c53"),
RAM_WORD'(x"8c170888"),
RAM_WORD'(x"1808718c"),
RAM_WORD'(x"120c8812"),
RAM_WORD'(x"0c587d51"),
RAM_WORD'(x"81f53f88"),
RAM_WORD'(x"1754f5bd"),
RAM_WORD'(x"39728415"),
RAM_WORD'(x"0cf41af8"),
RAM_WORD'(x"0670841e"),
RAM_WORD'(x"08810607"),
RAM_WORD'(x"841e0c70"),
RAM_WORD'(x"1d545b85"),
RAM_WORD'(x"0b84140c"),
RAM_WORD'(x"850b8814"),
RAM_WORD'(x"0c8f7b27"),
RAM_WORD'(x"fdcd3888"),
RAM_WORD'(x"1c527d51"),
RAM_WORD'(x"84d93f81"),
RAM_WORD'(x"87ec0b88"),
RAM_WORD'(x"05088187"),
RAM_WORD'(x"b0085955"),
RAM_WORD'(x"fdb53977"),
RAM_WORD'(x"8187b00c"),
RAM_WORD'(x"738187e0"),
RAM_WORD'(x"0cfc8939"),
RAM_WORD'(x"7284150c"),
RAM_WORD'(x"fda139f0"),
RAM_WORD'(x"3d0d7670"),
RAM_WORD'(x"797b5555"),
RAM_WORD'(x"55558f72"),
RAM_WORD'(x"278c3872"),
RAM_WORD'(x"75078306"),
RAM_WORD'(x"5170802e"),
RAM_WORD'(x"a938ff12"),
RAM_WORD'(x"5271ff2e"),
RAM_WORD'(x"98387270"),
RAM_WORD'(x"81055433"),
RAM_WORD'(x"74708105"),
RAM_WORD'(x"5634ff12"),
RAM_WORD'(x"5271ff2e"),
RAM_WORD'(x"098106ea"),
RAM_WORD'(x"38748190"),
RAM_WORD'(x"980c983d"),
RAM_WORD'(x"0d047451"),
RAM_WORD'(x"72708405"),
RAM_WORD'(x"54087170"),
RAM_WORD'(x"8405530c"),
RAM_WORD'(x"72708405"),
RAM_WORD'(x"54087170"),
RAM_WORD'(x"8405530c"),
RAM_WORD'(x"72708405"),
RAM_WORD'(x"54087170"),
RAM_WORD'(x"8405530c"),
RAM_WORD'(x"72708405"),
RAM_WORD'(x"54087170"),
RAM_WORD'(x"8405530c"),
RAM_WORD'(x"f0125271"),
RAM_WORD'(x"8f26c938"),
RAM_WORD'(x"83722795"),
RAM_WORD'(x"38727084"),
RAM_WORD'(x"05540871"),
RAM_WORD'(x"70840553"),
RAM_WORD'(x"0cfc1252"),
RAM_WORD'(x"718326ed"),
RAM_WORD'(x"387054ff"),
RAM_WORD'(x"81390404"),
RAM_WORD'(x"f43d0d80"),
RAM_WORD'(x"0b81e0a0"),
RAM_WORD'(x"0c7651eb"),
RAM_WORD'(x"d33f8190"),
RAM_WORD'(x"98085381"),
RAM_WORD'(x"909808ff"),
RAM_WORD'(x"2e8a3872"),
RAM_WORD'(x"8190980c"),
RAM_WORD'(x"943d0d04"),
RAM_WORD'(x"81e0a008"),
RAM_WORD'(x"5473802e"),
RAM_WORD'(x"ee387574"),
RAM_WORD'(x"710c5272"),
RAM_WORD'(x"8190980c"),
RAM_WORD'(x"943d0d04"),
RAM_WORD'(x"ec3d0d77"),
RAM_WORD'(x"79707207"),
RAM_WORD'(x"83065354"),
RAM_WORD'(x"52709338"),
RAM_WORD'(x"71737308"),
RAM_WORD'(x"54565471"),
RAM_WORD'(x"73082e80"),
RAM_WORD'(x"c6387375"),
RAM_WORD'(x"54527133"),
RAM_WORD'(x"7081ff06"),
RAM_WORD'(x"52547080"),
RAM_WORD'(x"2e9d3872"),
RAM_WORD'(x"33557075"),
RAM_WORD'(x"2e098106"),
RAM_WORD'(x"95388112"),
RAM_WORD'(x"81147133"),
RAM_WORD'(x"7081ff06"),
RAM_WORD'(x"54565452"),
RAM_WORD'(x"70e53872"),
RAM_WORD'(x"33557381"),
RAM_WORD'(x"ff067581"),
RAM_WORD'(x"ff067171"),
RAM_WORD'(x"31819098"),
RAM_WORD'(x"0c52529c"),
RAM_WORD'(x"3d0d0471"),
RAM_WORD'(x"0970f7fb"),
RAM_WORD'(x"fdff1406"),
RAM_WORD'(x"70f88482"),
RAM_WORD'(x"81800651"),
RAM_WORD'(x"51517097"),
RAM_WORD'(x"38841484"),
RAM_WORD'(x"16710854"),
RAM_WORD'(x"56547175"),
RAM_WORD'(x"082edc38"),
RAM_WORD'(x"73755452"),
RAM_WORD'(x"ff943980"),
RAM_WORD'(x"0b819098"),
RAM_WORD'(x"0c9c3d0d"),
RAM_WORD'(x"04ec3d0d"),
RAM_WORD'(x"77705256"),
RAM_WORD'(x"fea03f81"),
RAM_WORD'(x"87ec0b88"),
RAM_WORD'(x"05088411"),
RAM_WORD'(x"08fc0670"),
RAM_WORD'(x"7b319fef"),
RAM_WORD'(x"05e08006"),
RAM_WORD'(x"e0800556"),
RAM_WORD'(x"5653a080"),
RAM_WORD'(x"74249638"),
RAM_WORD'(x"80527551"),
RAM_WORD'(x"fdfa3f81"),
RAM_WORD'(x"87f40815"),
RAM_WORD'(x"53728190"),
RAM_WORD'(x"98082e91"),
RAM_WORD'(x"387551fd"),
RAM_WORD'(x"e63f8053"),
RAM_WORD'(x"72819098"),
RAM_WORD'(x"0c9c3d0d"),
RAM_WORD'(x"04733052"),
RAM_WORD'(x"7551fdd4"),
RAM_WORD'(x"3f819098"),
RAM_WORD'(x"08ff2eaa"),
RAM_WORD'(x"388187ec"),
RAM_WORD'(x"0b880508"),
RAM_WORD'(x"75753181"),
RAM_WORD'(x"0784120c"),
RAM_WORD'(x"538187b0"),
RAM_WORD'(x"08743181"),
RAM_WORD'(x"87b00c75"),
RAM_WORD'(x"51fdac3f"),
RAM_WORD'(x"810b8190"),
RAM_WORD'(x"980c9c3d"),
RAM_WORD'(x"0d048052"),
RAM_WORD'(x"7551fd9c"),
RAM_WORD'(x"3f8187ec"),
RAM_WORD'(x"0b880508"),
RAM_WORD'(x"81909808"),
RAM_WORD'(x"71315653"),
RAM_WORD'(x"8f7525ff"),
RAM_WORD'(x"9c388190"),
RAM_WORD'(x"98088187"),
RAM_WORD'(x"e0083181"),
RAM_WORD'(x"87b00c74"),
RAM_WORD'(x"81078414"),
RAM_WORD'(x"0c7551fc"),
RAM_WORD'(x"ee3f8053"),
RAM_WORD'(x"ff8639d8"),
RAM_WORD'(x"3d0d7c7e"),
RAM_WORD'(x"545b7280"),
RAM_WORD'(x"2e828338"),
RAM_WORD'(x"7a51fcd6"),
RAM_WORD'(x"3ff81384"),
RAM_WORD'(x"110870fe"),
RAM_WORD'(x"06701384"),
RAM_WORD'(x"1108fc06"),
RAM_WORD'(x"5d585954"),
RAM_WORD'(x"588187f4"),
RAM_WORD'(x"08752e82"),
RAM_WORD'(x"de387884"),
RAM_WORD'(x"160c8073"),
RAM_WORD'(x"8106545a"),
RAM_WORD'(x"727a2e81"),
RAM_WORD'(x"d5387815"),
RAM_WORD'(x"84110881"),
RAM_WORD'(x"06515372"),
RAM_WORD'(x"a0387817"),
RAM_WORD'(x"577981e6"),
RAM_WORD'(x"38881508"),
RAM_WORD'(x"53728187"),
RAM_WORD'(x"f42e82f9"),
RAM_WORD'(x"388c1508"),
RAM_WORD'(x"708c150c"),
RAM_WORD'(x"7388120c"),
RAM_WORD'(x"56768107"),
RAM_WORD'(x"84190c76"),
RAM_WORD'(x"1877710c"),
RAM_WORD'(x"53798191"),
RAM_WORD'(x"3883ff77"),
RAM_WORD'(x"2781c838"),
RAM_WORD'(x"76892a77"),
RAM_WORD'(x"832a5653"),
RAM_WORD'(x"72802ebf"),
RAM_WORD'(x"3876862a"),
RAM_WORD'(x"b8055584"),
RAM_WORD'(x"7327b438"),
RAM_WORD'(x"80db1355"),
RAM_WORD'(x"947327ab"),
RAM_WORD'(x"38768c2a"),
RAM_WORD'(x"80ee0555"),
RAM_WORD'(x"80d47327"),
RAM_WORD'(x"9e38768f"),
RAM_WORD'(x"2a80f705"),
RAM_WORD'(x"5582d473"),
RAM_WORD'(x"27913876"),
RAM_WORD'(x"922a80fc"),
RAM_WORD'(x"05558ad4"),
RAM_WORD'(x"73278438"),
RAM_WORD'(x"80fe5574"),
RAM_WORD'(x"10101081"),
RAM_WORD'(x"87ec0588"),
RAM_WORD'(x"11085556"),
RAM_WORD'(x"73762e82"),
RAM_WORD'(x"b3388414"),
RAM_WORD'(x"08fc0653"),
RAM_WORD'(x"7673278d"),
RAM_WORD'(x"38881408"),
RAM_WORD'(x"5473762e"),
RAM_WORD'(x"098106ea"),
RAM_WORD'(x"388c1408"),
RAM_WORD'(x"708c1a0c"),
RAM_WORD'(x"74881a0c"),
RAM_WORD'(x"7888120c"),
RAM_WORD'(x"56778c15"),
RAM_WORD'(x"0c7a51fa"),
RAM_WORD'(x"da3fb03d"),
RAM_WORD'(x"0d047708"),
RAM_WORD'(x"78713159"),
RAM_WORD'(x"77058819"),
RAM_WORD'(x"08545772"),
RAM_WORD'(x"8187f42e"),
RAM_WORD'(x"80e0388c"),
RAM_WORD'(x"1808708c"),
RAM_WORD'(x"150c7388"),
RAM_WORD'(x"120c56fe"),
RAM_WORD'(x"89398815"),
RAM_WORD'(x"088c1608"),
RAM_WORD'(x"708c130c"),
RAM_WORD'(x"5788170c"),
RAM_WORD'(x"fea33976"),
RAM_WORD'(x"832a7054"),
RAM_WORD'(x"55807524"),
RAM_WORD'(x"81983872"),
RAM_WORD'(x"822c8171"),
RAM_WORD'(x"2b8187f0"),
RAM_WORD'(x"08078187"),
RAM_WORD'(x"ec0b8405"),
RAM_WORD'(x"0c537410"),
RAM_WORD'(x"10108187"),
RAM_WORD'(x"ec058811"),
RAM_WORD'(x"08555675"),
RAM_WORD'(x"8c190c73"),
RAM_WORD'(x"88190c77"),
RAM_WORD'(x"88170c77"),
RAM_WORD'(x"8c150cff"),
RAM_WORD'(x"8439815a"),
RAM_WORD'(x"fdb43978"),
RAM_WORD'(x"17738106"),
RAM_WORD'(x"54577298"),
RAM_WORD'(x"38770878"),
RAM_WORD'(x"71315977"),
RAM_WORD'(x"058c1908"),
RAM_WORD'(x"881a0871"),
RAM_WORD'(x"8c120c88"),
RAM_WORD'(x"120c5757"),
RAM_WORD'(x"76810784"),
RAM_WORD'(x"190c7781"),
RAM_WORD'(x"87ec0b88"),
RAM_WORD'(x"050c8187"),
RAM_WORD'(x"e8087726"),
RAM_WORD'(x"fec73881"),
RAM_WORD'(x"87e40852"),
RAM_WORD'(x"7a51faf1"),
RAM_WORD'(x"3f7a51f9"),
RAM_WORD'(x"963ffeba"),
RAM_WORD'(x"3981788c"),
RAM_WORD'(x"150c7888"),
RAM_WORD'(x"150c738c"),
RAM_WORD'(x"1a0c7388"),
RAM_WORD'(x"1a0c5afd"),
RAM_WORD'(x"80398315"),
RAM_WORD'(x"70822c81"),
RAM_WORD'(x"712b8187"),
RAM_WORD'(x"f0080781"),
RAM_WORD'(x"87ec0b84"),
RAM_WORD'(x"050c5153"),
RAM_WORD'(x"74101010"),
RAM_WORD'(x"8187ec05"),
RAM_WORD'(x"88110855"),
RAM_WORD'(x"56fee439"),
RAM_WORD'(x"74538075"),
RAM_WORD'(x"24a73872"),
RAM_WORD'(x"822c8171"),
RAM_WORD'(x"2b8187f0"),
RAM_WORD'(x"08078187"),
RAM_WORD'(x"ec0b8405"),
RAM_WORD'(x"0c53758c"),
RAM_WORD'(x"190c7388"),
RAM_WORD'(x"190c7788"),
RAM_WORD'(x"170c778c"),
RAM_WORD'(x"150cfdcd"),
RAM_WORD'(x"39831570"),
RAM_WORD'(x"822c8171"),
RAM_WORD'(x"2b8187f0"),
RAM_WORD'(x"08078187"),
RAM_WORD'(x"ec0b8405"),
RAM_WORD'(x"0c5153d6"),
RAM_WORD'(x"3900ff39"),
RAM_WORD'(x"00ff39fc"),
RAM_WORD'(x"3d0d80d0"),
RAM_WORD'(x"ec0bfc05"),
RAM_WORD'(x"70085252"),
RAM_WORD'(x"70ff2e91"),
RAM_WORD'(x"38702dfc"),
RAM_WORD'(x"12700852"),
RAM_WORD'(x"5270ff2e"),
RAM_WORD'(x"098106f1"),
RAM_WORD'(x"388c3d0d"),
RAM_WORD'(x"0404d2fb"),
RAM_WORD'(x"3f040000"),
RAM_WORD'(x"00000001"),
RAM_WORD'(x"00000032"),
RAM_WORD'(x"64756d6d"),
RAM_WORD'(x"792e6578"),
RAM_WORD'(x"65000000"),
RAM_WORD'(x"30313233"),
RAM_WORD'(x"34353637"),
RAM_WORD'(x"38390000"),
RAM_WORD'(x"44485259"),
RAM_WORD'(x"53544f4e"),
RAM_WORD'(x"45205052"),
RAM_WORD'(x"4f475241"),
RAM_WORD'(x"4d2c2053"),
RAM_WORD'(x"4f4d4520"),
RAM_WORD'(x"53545249"),
RAM_WORD'(x"4e470000"),
RAM_WORD'(x"44485259"),
RAM_WORD'(x"53544f4e"),
RAM_WORD'(x"45205052"),
RAM_WORD'(x"4f475241"),
RAM_WORD'(x"4d2c2031"),
RAM_WORD'(x"27535420"),
RAM_WORD'(x"53545249"),
RAM_WORD'(x"4e470000"),
RAM_WORD'(x"44687279"),
RAM_WORD'(x"73746f6e"),
RAM_WORD'(x"65204265"),
RAM_WORD'(x"6e63686d"),
RAM_WORD'(x"61726b2c"),
RAM_WORD'(x"20566572"),
RAM_WORD'(x"73696f6e"),
RAM_WORD'(x"20322e31"),
RAM_WORD'(x"20284c61"),
RAM_WORD'(x"6e677561"),
RAM_WORD'(x"67653a20"),
RAM_WORD'(x"43290a00"),
RAM_WORD'(x"45786563"),
RAM_WORD'(x"7574696f"),
RAM_WORD'(x"6e207374"),
RAM_WORD'(x"61727473"),
RAM_WORD'(x"2c202564"),
RAM_WORD'(x"2072756e"),
RAM_WORD'(x"73207468"),
RAM_WORD'(x"726f7567"),
RAM_WORD'(x"68204468"),
RAM_WORD'(x"72797374"),
RAM_WORD'(x"6f6e650a"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"44485259"),
RAM_WORD'(x"53544f4e"),
RAM_WORD'(x"45205052"),
RAM_WORD'(x"4f475241"),
RAM_WORD'(x"4d2c2032"),
RAM_WORD'(x"274e4420"),
RAM_WORD'(x"53545249"),
RAM_WORD'(x"4e470000"),
RAM_WORD'(x"456e6420"),
RAM_WORD'(x"74696d65"),
RAM_WORD'(x"3a202564"),
RAM_WORD'(x"0a000000"),
RAM_WORD'(x"53746172"),
RAM_WORD'(x"74207469"),
RAM_WORD'(x"6d653a20"),
RAM_WORD'(x"25640a00"),
RAM_WORD'(x"45786563"),
RAM_WORD'(x"7574696f"),
RAM_WORD'(x"6e20656e"),
RAM_WORD'(x"64730a00"),
RAM_WORD'(x"75732f44"),
RAM_WORD'(x"68727973"),
RAM_WORD'(x"746f6e65"),
RAM_WORD'(x"3a200000"),
RAM_WORD'(x"44687279"),
RAM_WORD'(x"73746f6e"),
RAM_WORD'(x"652f7320"),
RAM_WORD'(x"3a200000"),
RAM_WORD'(x"2564200a"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"4d495053"),
RAM_WORD'(x"202a2031"),
RAM_WORD'(x"30303020"),
RAM_WORD'(x"3d202564"),
RAM_WORD'(x"200a0000"),
RAM_WORD'(x"46696e61"),
RAM_WORD'(x"6c207661"),
RAM_WORD'(x"6c756573"),
RAM_WORD'(x"206f6620"),
RAM_WORD'(x"74686520"),
RAM_WORD'(x"76617269"),
RAM_WORD'(x"61626c65"),
RAM_WORD'(x"73207573"),
RAM_WORD'(x"65642069"),
RAM_WORD'(x"6e207468"),
RAM_WORD'(x"65206265"),
RAM_WORD'(x"6e63686d"),
RAM_WORD'(x"61726b3a"),
RAM_WORD'(x"0a000000"),
RAM_WORD'(x"496e745f"),
RAM_WORD'(x"476c6f62"),
RAM_WORD'(x"3a202020"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"2025640a"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"73686f75"),
RAM_WORD'(x"6c642062"),
RAM_WORD'(x"653a2020"),
RAM_WORD'(x"2025640a"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"426f6f6c"),
RAM_WORD'(x"5f476c6f"),
RAM_WORD'(x"623a2020"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"2025640a"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"43685f31"),
RAM_WORD'(x"5f476c6f"),
RAM_WORD'(x"623a2020"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"2025630a"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"73686f75"),
RAM_WORD'(x"6c642062"),
RAM_WORD'(x"653a2020"),
RAM_WORD'(x"2025630a"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"43685f32"),
RAM_WORD'(x"5f476c6f"),
RAM_WORD'(x"623a2020"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"2025630a"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"4172725f"),
RAM_WORD'(x"315f476c"),
RAM_WORD'(x"6f625b38"),
RAM_WORD'(x"5d3a2020"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"2025640a"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"4172725f"),
RAM_WORD'(x"325f476c"),
RAM_WORD'(x"6f625b38"),
RAM_WORD'(x"5d5b375d"),
RAM_WORD'(x"3a202020"),
RAM_WORD'(x"2025640a"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"73686f75"),
RAM_WORD'(x"6c642062"),
RAM_WORD'(x"653a2020"),
RAM_WORD'(x"204e756d"),
RAM_WORD'(x"6265725f"),
RAM_WORD'(x"4f665f52"),
RAM_WORD'(x"756e7320"),
RAM_WORD'(x"2b203130"),
RAM_WORD'(x"0a000000"),
RAM_WORD'(x"5074725f"),
RAM_WORD'(x"476c6f62"),
RAM_WORD'(x"2d3e0a00"),
RAM_WORD'(x"20205074"),
RAM_WORD'(x"725f436f"),
RAM_WORD'(x"6d703a20"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"2025640a"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"73686f75"),
RAM_WORD'(x"6c642062"),
RAM_WORD'(x"653a2020"),
RAM_WORD'(x"2028696d"),
RAM_WORD'(x"706c656d"),
RAM_WORD'(x"656e7461"),
RAM_WORD'(x"74696f6e"),
RAM_WORD'(x"2d646570"),
RAM_WORD'(x"656e6465"),
RAM_WORD'(x"6e74290a"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"20204469"),
RAM_WORD'(x"7363723a"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"2025640a"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"2020456e"),
RAM_WORD'(x"756d5f43"),
RAM_WORD'(x"6f6d703a"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"2025640a"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"2020496e"),
RAM_WORD'(x"745f436f"),
RAM_WORD'(x"6d703a20"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"2025640a"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"20205374"),
RAM_WORD'(x"725f436f"),
RAM_WORD'(x"6d703a20"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"2025730a"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"73686f75"),
RAM_WORD'(x"6c642062"),
RAM_WORD'(x"653a2020"),
RAM_WORD'(x"20444852"),
RAM_WORD'(x"5953544f"),
RAM_WORD'(x"4e452050"),
RAM_WORD'(x"524f4752"),
RAM_WORD'(x"414d2c20"),
RAM_WORD'(x"534f4d45"),
RAM_WORD'(x"20535452"),
RAM_WORD'(x"494e470a"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"4e657874"),
RAM_WORD'(x"5f507472"),
RAM_WORD'(x"5f476c6f"),
RAM_WORD'(x"622d3e0a"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"73686f75"),
RAM_WORD'(x"6c642062"),
RAM_WORD'(x"653a2020"),
RAM_WORD'(x"2028696d"),
RAM_WORD'(x"706c656d"),
RAM_WORD'(x"656e7461"),
RAM_WORD'(x"74696f6e"),
RAM_WORD'(x"2d646570"),
RAM_WORD'(x"656e6465"),
RAM_WORD'(x"6e74292c"),
RAM_WORD'(x"2073616d"),
RAM_WORD'(x"65206173"),
RAM_WORD'(x"2061626f"),
RAM_WORD'(x"76650a00"),
RAM_WORD'(x"496e745f"),
RAM_WORD'(x"315f4c6f"),
RAM_WORD'(x"633a2020"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"2025640a"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"496e745f"),
RAM_WORD'(x"325f4c6f"),
RAM_WORD'(x"633a2020"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"2025640a"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"496e745f"),
RAM_WORD'(x"335f4c6f"),
RAM_WORD'(x"633a2020"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"2025640a"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"456e756d"),
RAM_WORD'(x"5f4c6f63"),
RAM_WORD'(x"3a202020"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"2025640a"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"5374725f"),
RAM_WORD'(x"315f4c6f"),
RAM_WORD'(x"633a2020"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"2025730a"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"73686f75"),
RAM_WORD'(x"6c642062"),
RAM_WORD'(x"653a2020"),
RAM_WORD'(x"20444852"),
RAM_WORD'(x"5953544f"),
RAM_WORD'(x"4e452050"),
RAM_WORD'(x"524f4752"),
RAM_WORD'(x"414d2c20"),
RAM_WORD'(x"31275354"),
RAM_WORD'(x"20535452"),
RAM_WORD'(x"494e470a"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"5374725f"),
RAM_WORD'(x"325f4c6f"),
RAM_WORD'(x"633a2020"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"2025730a"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"20202020"),
RAM_WORD'(x"73686f75"),
RAM_WORD'(x"6c642062"),
RAM_WORD'(x"653a2020"),
RAM_WORD'(x"20444852"),
RAM_WORD'(x"5953544f"),
RAM_WORD'(x"4e452050"),
RAM_WORD'(x"524f4752"),
RAM_WORD'(x"414d2c20"),
RAM_WORD'(x"32274e44"),
RAM_WORD'(x"20535452"),
RAM_WORD'(x"494e470a"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"44485259"),
RAM_WORD'(x"53544f4e"),
RAM_WORD'(x"45205052"),
RAM_WORD'(x"4f475241"),
RAM_WORD'(x"4d2c2033"),
RAM_WORD'(x"27524420"),
RAM_WORD'(x"53545249"),
RAM_WORD'(x"4e470000"),
RAM_WORD'(x"43000000"),
RAM_WORD'(x"00ffffff"),
RAM_WORD'(x"ff00ffff"),
RAM_WORD'(x"ffff00ff"),
RAM_WORD'(x"ffffff00"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00002874"),
RAM_WORD'(x"0000c000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00007024"),
RAM_WORD'(x"00001b58"),
RAM_WORD'(x"00004034"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"0000429c"),
RAM_WORD'(x"000042f8"),
RAM_WORD'(x"00004354"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00002070"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000001"),
RAM_WORD'(x"330eabcd"),
RAM_WORD'(x"1234e66d"),
RAM_WORD'(x"deec0005"),
RAM_WORD'(x"000b0000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"ffffffff"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00020000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"000043ec"),
RAM_WORD'(x"000043ec"),
RAM_WORD'(x"000043f4"),
RAM_WORD'(x"000043f4"),
RAM_WORD'(x"000043fc"),
RAM_WORD'(x"000043fc"),
RAM_WORD'(x"00004404"),
RAM_WORD'(x"00004404"),
RAM_WORD'(x"0000440c"),
RAM_WORD'(x"0000440c"),
RAM_WORD'(x"00004414"),
RAM_WORD'(x"00004414"),
RAM_WORD'(x"0000441c"),
RAM_WORD'(x"0000441c"),
RAM_WORD'(x"00004424"),
RAM_WORD'(x"00004424"),
RAM_WORD'(x"0000442c"),
RAM_WORD'(x"0000442c"),
RAM_WORD'(x"00004434"),
RAM_WORD'(x"00004434"),
RAM_WORD'(x"0000443c"),
RAM_WORD'(x"0000443c"),
RAM_WORD'(x"00004444"),
RAM_WORD'(x"00004444"),
RAM_WORD'(x"0000444c"),
RAM_WORD'(x"0000444c"),
RAM_WORD'(x"00004454"),
RAM_WORD'(x"00004454"),
RAM_WORD'(x"0000445c"),
RAM_WORD'(x"0000445c"),
RAM_WORD'(x"00004464"),
RAM_WORD'(x"00004464"),
RAM_WORD'(x"0000446c"),
RAM_WORD'(x"0000446c"),
RAM_WORD'(x"00004474"),
RAM_WORD'(x"00004474"),
RAM_WORD'(x"0000447c"),
RAM_WORD'(x"0000447c"),
RAM_WORD'(x"00004484"),
RAM_WORD'(x"00004484"),
RAM_WORD'(x"0000448c"),
RAM_WORD'(x"0000448c"),
RAM_WORD'(x"00004494"),
RAM_WORD'(x"00004494"),
RAM_WORD'(x"0000449c"),
RAM_WORD'(x"0000449c"),
RAM_WORD'(x"000044a4"),
RAM_WORD'(x"000044a4"),
RAM_WORD'(x"000044ac"),
RAM_WORD'(x"000044ac"),
RAM_WORD'(x"000044b4"),
RAM_WORD'(x"000044b4"),
RAM_WORD'(x"000044bc"),
RAM_WORD'(x"000044bc"),
RAM_WORD'(x"000044c4"),
RAM_WORD'(x"000044c4"),
RAM_WORD'(x"000044cc"),
RAM_WORD'(x"000044cc"),
RAM_WORD'(x"000044d4"),
RAM_WORD'(x"000044d4"),
RAM_WORD'(x"000044dc"),
RAM_WORD'(x"000044dc"),
RAM_WORD'(x"000044e4"),
RAM_WORD'(x"000044e4"),
RAM_WORD'(x"000044ec"),
RAM_WORD'(x"000044ec"),
RAM_WORD'(x"000044f4"),
RAM_WORD'(x"000044f4"),
RAM_WORD'(x"000044fc"),
RAM_WORD'(x"000044fc"),
RAM_WORD'(x"00004504"),
RAM_WORD'(x"00004504"),
RAM_WORD'(x"0000450c"),
RAM_WORD'(x"0000450c"),
RAM_WORD'(x"00004514"),
RAM_WORD'(x"00004514"),
RAM_WORD'(x"0000451c"),
RAM_WORD'(x"0000451c"),
RAM_WORD'(x"00004524"),
RAM_WORD'(x"00004524"),
RAM_WORD'(x"0000452c"),
RAM_WORD'(x"0000452c"),
RAM_WORD'(x"00004534"),
RAM_WORD'(x"00004534"),
RAM_WORD'(x"0000453c"),
RAM_WORD'(x"0000453c"),
RAM_WORD'(x"00004544"),
RAM_WORD'(x"00004544"),
RAM_WORD'(x"0000454c"),
RAM_WORD'(x"0000454c"),
RAM_WORD'(x"00004554"),
RAM_WORD'(x"00004554"),
RAM_WORD'(x"0000455c"),
RAM_WORD'(x"0000455c"),
RAM_WORD'(x"00004564"),
RAM_WORD'(x"00004564"),
RAM_WORD'(x"0000456c"),
RAM_WORD'(x"0000456c"),
RAM_WORD'(x"00004574"),
RAM_WORD'(x"00004574"),
RAM_WORD'(x"0000457c"),
RAM_WORD'(x"0000457c"),
RAM_WORD'(x"00004584"),
RAM_WORD'(x"00004584"),
RAM_WORD'(x"0000458c"),
RAM_WORD'(x"0000458c"),
RAM_WORD'(x"00004594"),
RAM_WORD'(x"00004594"),
RAM_WORD'(x"0000459c"),
RAM_WORD'(x"0000459c"),
RAM_WORD'(x"000045a4"),
RAM_WORD'(x"000045a4"),
RAM_WORD'(x"000045ac"),
RAM_WORD'(x"000045ac"),
RAM_WORD'(x"000045b4"),
RAM_WORD'(x"000045b4"),
RAM_WORD'(x"000045bc"),
RAM_WORD'(x"000045bc"),
RAM_WORD'(x"000045c4"),
RAM_WORD'(x"000045c4"),
RAM_WORD'(x"000045cc"),
RAM_WORD'(x"000045cc"),
RAM_WORD'(x"000045d4"),
RAM_WORD'(x"000045d4"),
RAM_WORD'(x"000045dc"),
RAM_WORD'(x"000045dc"),
RAM_WORD'(x"000045e4"),
RAM_WORD'(x"000045e4"),
RAM_WORD'(x"000045ec"),
RAM_WORD'(x"000045ec"),
RAM_WORD'(x"000045f4"),
RAM_WORD'(x"000045f4"),
RAM_WORD'(x"000045fc"),
RAM_WORD'(x"000045fc"),
RAM_WORD'(x"00004604"),
RAM_WORD'(x"00004604"),
RAM_WORD'(x"0000460c"),
RAM_WORD'(x"0000460c"),
RAM_WORD'(x"00004614"),
RAM_WORD'(x"00004614"),
RAM_WORD'(x"0000461c"),
RAM_WORD'(x"0000461c"),
RAM_WORD'(x"00004624"),
RAM_WORD'(x"00004624"),
RAM_WORD'(x"0000462c"),
RAM_WORD'(x"0000462c"),
RAM_WORD'(x"00004634"),
RAM_WORD'(x"00004634"),
RAM_WORD'(x"0000463c"),
RAM_WORD'(x"0000463c"),
RAM_WORD'(x"00004644"),
RAM_WORD'(x"00004644"),
RAM_WORD'(x"0000464c"),
RAM_WORD'(x"0000464c"),
RAM_WORD'(x"00004654"),
RAM_WORD'(x"00004654"),
RAM_WORD'(x"0000465c"),
RAM_WORD'(x"0000465c"),
RAM_WORD'(x"00004664"),
RAM_WORD'(x"00004664"),
RAM_WORD'(x"0000466c"),
RAM_WORD'(x"0000466c"),
RAM_WORD'(x"00004674"),
RAM_WORD'(x"00004674"),
RAM_WORD'(x"0000467c"),
RAM_WORD'(x"0000467c"),
RAM_WORD'(x"00004684"),
RAM_WORD'(x"00004684"),
RAM_WORD'(x"0000468c"),
RAM_WORD'(x"0000468c"),
RAM_WORD'(x"00004694"),
RAM_WORD'(x"00004694"),
RAM_WORD'(x"0000469c"),
RAM_WORD'(x"0000469c"),
RAM_WORD'(x"000046a4"),
RAM_WORD'(x"000046a4"),
RAM_WORD'(x"000046ac"),
RAM_WORD'(x"000046ac"),
RAM_WORD'(x"000046b4"),
RAM_WORD'(x"000046b4"),
RAM_WORD'(x"000046bc"),
RAM_WORD'(x"000046bc"),
RAM_WORD'(x"000046c4"),
RAM_WORD'(x"000046c4"),
RAM_WORD'(x"000046cc"),
RAM_WORD'(x"000046cc"),
RAM_WORD'(x"000046d4"),
RAM_WORD'(x"000046d4"),
RAM_WORD'(x"000046dc"),
RAM_WORD'(x"000046dc"),
RAM_WORD'(x"000046e4"),
RAM_WORD'(x"000046e4"),
RAM_WORD'(x"000046ec"),
RAM_WORD'(x"000046ec"),
RAM_WORD'(x"000046f4"),
RAM_WORD'(x"000046f4"),
RAM_WORD'(x"000046fc"),
RAM_WORD'(x"000046fc"),
RAM_WORD'(x"00004704"),
RAM_WORD'(x"00004704"),
RAM_WORD'(x"0000470c"),
RAM_WORD'(x"0000470c"),
RAM_WORD'(x"00004714"),
RAM_WORD'(x"00004714"),
RAM_WORD'(x"0000471c"),
RAM_WORD'(x"0000471c"),
RAM_WORD'(x"00004724"),
RAM_WORD'(x"00004724"),
RAM_WORD'(x"0000472c"),
RAM_WORD'(x"0000472c"),
RAM_WORD'(x"00004734"),
RAM_WORD'(x"00004734"),
RAM_WORD'(x"0000473c"),
RAM_WORD'(x"0000473c"),
RAM_WORD'(x"00004744"),
RAM_WORD'(x"00004744"),
RAM_WORD'(x"0000474c"),
RAM_WORD'(x"0000474c"),
RAM_WORD'(x"00004754"),
RAM_WORD'(x"00004754"),
RAM_WORD'(x"0000475c"),
RAM_WORD'(x"0000475c"),
RAM_WORD'(x"00004764"),
RAM_WORD'(x"00004764"),
RAM_WORD'(x"0000476c"),
RAM_WORD'(x"0000476c"),
RAM_WORD'(x"00004774"),
RAM_WORD'(x"00004774"),
RAM_WORD'(x"0000477c"),
RAM_WORD'(x"0000477c"),
RAM_WORD'(x"00004784"),
RAM_WORD'(x"00004784"),
RAM_WORD'(x"0000478c"),
RAM_WORD'(x"0000478c"),
RAM_WORD'(x"00004794"),
RAM_WORD'(x"00004794"),
RAM_WORD'(x"0000479c"),
RAM_WORD'(x"0000479c"),
RAM_WORD'(x"000047a4"),
RAM_WORD'(x"000047a4"),
RAM_WORD'(x"000047ac"),
RAM_WORD'(x"000047ac"),
RAM_WORD'(x"000047b4"),
RAM_WORD'(x"000047b4"),
RAM_WORD'(x"000047bc"),
RAM_WORD'(x"000047bc"),
RAM_WORD'(x"000047c4"),
RAM_WORD'(x"000047c4"),
RAM_WORD'(x"000047cc"),
RAM_WORD'(x"000047cc"),
RAM_WORD'(x"000047d4"),
RAM_WORD'(x"000047d4"),
RAM_WORD'(x"000047dc"),
RAM_WORD'(x"000047dc"),
RAM_WORD'(x"000047e4"),
RAM_WORD'(x"000047e4"),
RAM_WORD'(x"ffffffff"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"ffffffff"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000")
);

begin

  process (clk)
  begin
    if rising_edge(clk) then
      if memAWriteEnable='1' then
        RAM( conv_integer(memAAddr) ) := memAWrite;
      end if;
      memARead <= RAM(conv_integer(memAAddr)) ;
    end if;
  end process;  

  process (clk)
  begin
    if rising_edge(clk) then
      if memBWriteEnable='1' then
        RAM( conv_integer(memBAddr) ) := memBWrite;
      end if;
      memBRead <= RAM(conv_integer(memBAddr)) ;
    end if;
  end process;  

end behave; 
