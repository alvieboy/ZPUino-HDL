library IEEE; 
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
library UNISIM;
use UNISIM.vcomponents.all;
entity dp_rom_32_32 is 
port (ADDRA: in std_logic_vector(13 downto 2);
      CLK : in std_logic;
      ENA:   in std_logic;
      WEA: in std_logic; -- to avoid a bug in Xilinx ISE
      DOA: out STD_LOGIC_VECTOR (31 downto 0);
      ADDRB: in std_logic_vector(13 downto 2);
      DIA: in STD_LOGIC_VECTOR (31 downto 0); -- to avoid a bug in Xilinx ISE
      WEB: in std_logic;
      ENB:   in std_logic;
      DOB: out STD_LOGIC_VECTOR (31 downto 0);
      DIB: in STD_LOGIC_VECTOR (31 downto 0));
end dp_rom_32_32;
architecture behave of dp_rom_32_32 is
signal ram_0_DOB: std_logic_vector(3 downto 0);
signal ram_0_DIB: std_logic_vector(3 downto 0);
signal ram_0_DOA: std_logic_vector(3 downto 0);
signal ram_0_DIA: std_logic_vector(3 downto 0);
signal ram_1_DOB: std_logic_vector(3 downto 0);
signal ram_1_DIB: std_logic_vector(3 downto 0);
signal ram_1_DOA: std_logic_vector(3 downto 0);
signal ram_1_DIA: std_logic_vector(3 downto 0);
signal ram_2_DOB: std_logic_vector(3 downto 0);
signal ram_2_DIB: std_logic_vector(3 downto 0);
signal ram_2_DOA: std_logic_vector(3 downto 0);
signal ram_2_DIA: std_logic_vector(3 downto 0);
signal ram_3_DOB: std_logic_vector(3 downto 0);
signal ram_3_DIB: std_logic_vector(3 downto 0);
signal ram_3_DOA: std_logic_vector(3 downto 0);
signal ram_3_DIA: std_logic_vector(3 downto 0);
signal ram_4_DOB: std_logic_vector(3 downto 0);
signal ram_4_DIB: std_logic_vector(3 downto 0);
signal ram_4_DOA: std_logic_vector(3 downto 0);
signal ram_4_DIA: std_logic_vector(3 downto 0);
signal ram_5_DOB: std_logic_vector(3 downto 0);
signal ram_5_DIB: std_logic_vector(3 downto 0);
signal ram_5_DOA: std_logic_vector(3 downto 0);
signal ram_5_DIA: std_logic_vector(3 downto 0);
signal ram_6_DOB: std_logic_vector(3 downto 0);
signal ram_6_DIB: std_logic_vector(3 downto 0);
signal ram_6_DOA: std_logic_vector(3 downto 0);
signal ram_6_DIA: std_logic_vector(3 downto 0);
signal ram_7_DOB: std_logic_vector(3 downto 0);
signal ram_7_DIB: std_logic_vector(3 downto 0);
signal ram_7_DOA: std_logic_vector(3 downto 0);
signal ram_7_DIA: std_logic_vector(3 downto 0);

begin
DOB(0) <= ram_0_DOB(3);
DOB(1) <= ram_1_DOB(3);
DOB(2) <= ram_2_DOB(3);
DOB(3) <= ram_3_DOB(3);
DOB(4) <= ram_4_DOB(3);
DOB(5) <= ram_5_DOB(3);
DOB(6) <= ram_6_DOB(3);
DOB(7) <= ram_7_DOB(3);
DOB(8) <= ram_0_DOB(2);
DOB(9) <= ram_1_DOB(2);
DOB(10) <= ram_2_DOB(2);
DOB(11) <= ram_3_DOB(2);
DOB(12) <= ram_4_DOB(2);
DOB(13) <= ram_5_DOB(2);
DOB(14) <= ram_6_DOB(2);
DOB(15) <= ram_7_DOB(2);
DOB(16) <= ram_0_DOB(1);
DOB(17) <= ram_1_DOB(1);
DOB(18) <= ram_2_DOB(1);
DOB(19) <= ram_3_DOB(1);
DOB(20) <= ram_4_DOB(1);
DOB(21) <= ram_5_DOB(1);
DOB(22) <= ram_6_DOB(1);
DOB(23) <= ram_7_DOB(1);
DOB(24) <= ram_0_DOB(0);
DOB(25) <= ram_1_DOB(0);
DOB(26) <= ram_2_DOB(0);
DOB(27) <= ram_3_DOB(0);
DOB(28) <= ram_4_DOB(0);
DOB(29) <= ram_5_DOB(0);
DOB(30) <= ram_6_DOB(0);
DOB(31) <= ram_7_DOB(0);
DOA(0) <= ram_0_DOA(3);
DOA(1) <= ram_1_DOA(3);
DOA(2) <= ram_2_DOA(3);
DOA(3) <= ram_3_DOA(3);
DOA(4) <= ram_4_DOA(3);
DOA(5) <= ram_5_DOA(3);
DOA(6) <= ram_6_DOA(3);
DOA(7) <= ram_7_DOA(3);
DOA(8) <= ram_0_DOA(2);
DOA(9) <= ram_1_DOA(2);
DOA(10) <= ram_2_DOA(2);
DOA(11) <= ram_3_DOA(2);
DOA(12) <= ram_4_DOA(2);
DOA(13) <= ram_5_DOA(2);
DOA(14) <= ram_6_DOA(2);
DOA(15) <= ram_7_DOA(2);
DOA(16) <= ram_0_DOA(1);
DOA(17) <= ram_1_DOA(1);
DOA(18) <= ram_2_DOA(1);
DOA(19) <= ram_3_DOA(1);
DOA(20) <= ram_4_DOA(1);
DOA(21) <= ram_5_DOA(1);
DOA(22) <= ram_6_DOA(1);
DOA(23) <= ram_7_DOA(1);
DOA(24) <= ram_0_DOA(0);
DOA(25) <= ram_1_DOA(0);
DOA(26) <= ram_2_DOA(0);
DOA(27) <= ram_3_DOA(0);
DOA(28) <= ram_4_DOA(0);
DOA(29) <= ram_5_DOA(0);
DOA(30) <= ram_6_DOA(0);
DOA(31) <= ram_7_DOA(0);
ram_0_DIA(3) <= DIA(0);
ram_1_DIA(3) <= DIA(1);
ram_2_DIA(3) <= DIA(2);
ram_3_DIA(3) <= DIA(3);
ram_4_DIA(3) <= DIA(4);
ram_5_DIA(3) <= DIA(5);
ram_6_DIA(3) <= DIA(6);
ram_7_DIA(3) <= DIA(7);
ram_0_DIA(2) <= DIA(8);
ram_1_DIA(2) <= DIA(9);
ram_2_DIA(2) <= DIA(10);
ram_3_DIA(2) <= DIA(11);
ram_4_DIA(2) <= DIA(12);
ram_5_DIA(2) <= DIA(13);
ram_6_DIA(2) <= DIA(14);
ram_7_DIA(2) <= DIA(15);
ram_0_DIA(1) <= DIA(16);
ram_1_DIA(1) <= DIA(17);
ram_2_DIA(1) <= DIA(18);
ram_3_DIA(1) <= DIA(19);
ram_4_DIA(1) <= DIA(20);
ram_5_DIA(1) <= DIA(21);
ram_6_DIA(1) <= DIA(22);
ram_7_DIA(1) <= DIA(23);
ram_0_DIA(0) <= DIA(24);
ram_1_DIA(0) <= DIA(25);
ram_2_DIA(0) <= DIA(26);
ram_3_DIA(0) <= DIA(27);
ram_4_DIA(0) <= DIA(28);
ram_5_DIA(0) <= DIA(29);
ram_6_DIA(0) <= DIA(30);
ram_7_DIA(0) <= DIA(31);
ram_0_DIB(3) <= DIB(0);
ram_1_DIB(3) <= DIB(1);
ram_2_DIB(3) <= DIB(2);
ram_3_DIB(3) <= DIB(3);
ram_4_DIB(3) <= DIB(4);
ram_5_DIB(3) <= DIB(5);
ram_6_DIB(3) <= DIB(6);
ram_7_DIB(3) <= DIB(7);
ram_0_DIB(2) <= DIB(8);
ram_1_DIB(2) <= DIB(9);
ram_2_DIB(2) <= DIB(10);
ram_3_DIB(2) <= DIB(11);
ram_4_DIB(2) <= DIB(12);
ram_5_DIB(2) <= DIB(13);
ram_6_DIB(2) <= DIB(14);
ram_7_DIB(2) <= DIB(15);
ram_0_DIB(1) <= DIB(16);
ram_1_DIB(1) <= DIB(17);
ram_2_DIB(1) <= DIB(18);
ram_3_DIB(1) <= DIB(19);
ram_4_DIB(1) <= DIB(20);
ram_5_DIB(1) <= DIB(21);
ram_6_DIB(1) <= DIB(22);
ram_7_DIB(1) <= DIB(23);
ram_0_DIB(0) <= DIB(24);
ram_1_DIB(0) <= DIB(25);
ram_2_DIB(0) <= DIB(26);
ram_3_DIB(0) <= DIB(27);
ram_4_DIB(0) <= DIB(28);
ram_5_DIB(0) <= DIB(29);
ram_6_DIB(0) <= DIB(30);
ram_7_DIB(0) <= DIB(31);
RAM_0_inst : RAMB16_S4_S4 
generic map ( 
INIT_00 => X"000001d803d6005f000001d8003575ee3ff7ddf30003bba30000000700000017",
INIT_01 => X"0003676e0001a76e061fbb2f000ed538000013f4000000680000001700000000",
INIT_02 => X"0f734d3a0000001700000017002e467100030fa100000772000000fc0000000f",
INIT_03 => X"000002ff000000000000004400000000000000070000011f000000071ee69b3a",
INIT_04 => X"de7659780f8e3e004000019f80c02003602002603d40ce80c31f6ec000000025",
INIT_05 => X"4d9ec7ad01f56fa4bc00f6d07f3666c1fb36b8d97bb0067ceb076dec05d20306",
INIT_06 => X"864cd1fd99c0020238004040404810080f4f8b14470300ee1001c381018e0718",
INIT_07 => X"309b0004078180bb359af9cab0009f77040cfcff0187aa043d52194001700002",
INIT_08 => X"e77b29c997cb8f800264e6ffd703d1f679bffddbe6560b6ffdf35e8ff19dffdf",
INIT_09 => X"6f677be9fedbffed67f00b00024f0080e07c9fc7003f02f03fcdff81f402d9ed",
INIT_0A => X"e31fe6b2793e43e49f8448606979f67ba93f3eed653f7a1f7d28742e7020da40",
INIT_0B => X"f8f8fbb0201006066b2d4af58c1a579e7fde79f9f1027bf0f9c1f696cd6c7d9a",
INIT_0C => X"3c9821f63f3c7c07c07a93e9f8d1c3e03c60403ca7c7d00b4d05023060540c18",
INIT_0D => X"000000000000000256141ccc44000087bde0875a025053bf8ec181401a1e3f1f",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"000000000000000000000000000000000000000000000000000000000f0f4000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000100",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map ( 
DOA => ram_0_DOA, -- 4-bit Data Output 
ADDRA => ADDRA, -- 14-bit Address Input 
CLKA => CLK, -- Clock 
DIA => ram_0_DIA, -- 4-bit Data Input 
ENA => ENA, -- RAM Enable Input 
WEA => WEA, -- Write Enable Input 
DOB => ram_0_DOB, -- 4-bit Data Output 
ADDRB => ADDRB, -- 12-bit Address Input 
CLKB => CLK, -- Clock 
SSRA => '0', 
SSRB => '0', 
DIB => ram_0_DIB, -- 4-bit Data Input 
ENB => ENB, -- RAM Enable Input 
WEB => WEB -- Write Enable Input 
);
RAM_1_inst : RAMB16_S4_S4 
generic map ( 
INIT_00 => X"000000ff012976a2000000fb001bdad13ffba3f4000ff4740000001f0000000f",
INIT_01 => X"000198110000d81100bf4794000768ff00000b8f0000003f0000001700000000",
INIT_02 => X"01a586c10000001700000017000f0ef4000e8474000003bd0000004300000010",
INIT_03 => X"00000148000000000000008900000000000000080000001e00000002034b0cc1",
INIT_04 => X"bcf1257b1e023c300266049c802000408000418010ee33581708fa400000003c",
INIT_05 => X"090e2382005042d161e291697c01ca137883556091e0010436b3cc02b4240001",
INIT_06 => X"8e4815f597c0020278004040404010080c02821441df0023b8004b8101e22952",
INIT_07 => X"084600040401882009296044c8388f11de2870722b92494a124d54e811f00002",
INIT_08 => X"8b79629521a30f40022d0affdf0212f762fef004e8381e7b7fe0df2fc047f7b0",
INIT_09 => X"34c9abedfe4fef024a680830558680c0e0405fd5302f02f03f17f78102030009",
INIT_0A => X"8b0f0024321ca1ca0e5148d00298f112cc431e204a535c0d1a5836090022a480",
INIT_0B => X"78787886c0199f01000836f2615a478e3b9e38e8ee037baafab8f10d02d03c05",
INIT_0C => X"1c6608f31c1d7b03cc39c1c8f12011e61c98531c63c3c8082096024240440c14",
INIT_0D => X"0000000000000001740404c08c484447bde0a126c836148b22292000008e1e5f",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"000000000000000000000000000000000000000000000000000000000f0f4000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000100",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map ( 
DOA => ram_1_DOA, -- 4-bit Data Output 
ADDRA => ADDRA, -- 14-bit Address Input 
CLKA => CLK, -- Clock 
DIA => ram_1_DIA, -- 4-bit Data Input 
ENA => ENA, -- RAM Enable Input 
WEA => WEA, -- Write Enable Input 
DOB => ram_1_DOB, -- 4-bit Data Output 
ADDRB => ADDRB, -- 12-bit Address Input 
CLKB => CLK, -- Clock 
SSRA => '0', 
SSRB => '0', 
DIB => ram_1_DIB, -- 4-bit Data Input 
ENB => ENB, -- RAM Enable Input 
WEB => WEB -- Write Enable Input 
);
RAM_2_inst : RAMB16_S4_S4 
generic map ( 
INIT_00 => X"00000264042400a00000026400498a2860c8526600170a460000002000000020",
INIT_01 => X"00048a2800024a2809d0a4e00013e2680000384c000000800000002000000000",
INIT_02 => X"11f8ae5000000030000000300041490600160a46000009880000013000000028",
INIT_03 => X"0000061c00000000000001460000000000000014000002c00000000f23f15c50",
INIT_04 => X"a08e640311bd800051200443eea2574362574362410067073a14990000000066",
INIT_05 => X"1930042225db5d9464007eca1b7a61831ffe00c984e44ff76630c3fd04204b7e",
INIT_06 => X"5df62864d790c0c0f21818181806030703cccaca0e2b10fc5021f0e444dd0684",
INIT_07 => X"f4e62181826098ff7688dba04909b07e2e03818fd38381609c8a0eb21d1890c0",
INIT_08 => X"200188408b706010c070c10011c18d0210000ffc3c8cb9868212200022000053",
INIT_09 => X"65462408040000ffa2df07bfa48ff030382ec4069c10c10c00800060bfc1fff2",
INIT_0A => X"b0506fd07862062070e29148783707ed9106e0ffa106041d4208763ffca48409",
INIT_0B => X"838283f962070687f8226002420c1011460045190088010c308107f4dd5f41ba",
INIT_0C => X"a0e60f01a22200140c41820d0330de0220985060d41c1f07ffe0c83c18172186",
INIT_0D => X"0000000000000000051448c808880087bde1be2606306ff70fd05d0099d0e086",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"000000000000000000000000000000000000000000000000000000000f0fc000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map ( 
DOA => ram_2_DOA, -- 4-bit Data Output 
ADDRA => ADDRA, -- 14-bit Address Input 
CLKA => CLK, -- Clock 
DIA => ram_2_DIA, -- 4-bit Data Input 
ENA => ENA, -- RAM Enable Input 
WEA => WEA, -- Write Enable Input 
DOB => ram_2_DOB, -- 4-bit Data Output 
ADDRB => ADDRB, -- 12-bit Address Input 
CLKB => CLK, -- Clock 
SSRA => '0', 
SSRB => '0', 
DIB => ram_2_DIB, -- 4-bit Data Input 
ENB => ENB, -- RAM Enable Input 
WEB => WEB -- Write Enable Input 
);
RAM_3_inst : RAMB16_S4_S4 
generic map ( 
INIT_00 => X"000000200009540800000020000225020fc7046a0003608a0000001f0000001f",
INIT_01 => X"0000344200001442014e082000004dac000007940000001a0000000f00000000",
INIT_02 => X"002204a20000001f0000000f003e80fa0002808a000000420000000400000002",
INIT_03 => X"0000020800000000000000000000000000000000000000de00000002004409a2",
INIT_04 => X"9cf68d7f5f8cbd0b58a1685fbeb79f32979f329783280a022901080000000024",
INIT_05 => X"325f9fc041f3cd57273676ab3b36780b0bb520ab00a64768527040ed8c048306",
INIT_06 => X"3c684cee11a08282341050505044160a0e8fae96462742ec4885d9c5658de7c6",
INIT_07 => X"b6e2410505c13bb737e0b9b119017f7626a2f2ffd9b74f493af8cf94021ca082",
INIT_08 => X"38fc0e76e2f81f2082c021f7f18001fc087dfbdb20005812ffe03e87d0c3eff7",
INIT_09 => X"55d007f0fb47dfedf8be0ac0083fe020306bc7e0081f81f81f43efc1af82bdbe",
INIT_0A => X"997f66fdfeffbffa7eea91405e2df76f59c5beedf9c581ffc017faef68018090",
INIT_0B => X"fafbfbb108442e17688cd1fcc0c30fdf7a3f7dedf8c8fc0e7405f7fdcdcbfd9b",
INIT_0C => X"bd4eeff7bcbcf87fddfc8bfff677efeebf3bd0ffbfdfde0afbf48bae50720896",
INIT_0D => X"000000000000000004642c84c4c44c47bde0a68e26b137b40ed97d25fafefece",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"000000000000000000000000000000000000000000000000000000000f0fc000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000100",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map ( 
DOA => ram_3_DOA, -- 4-bit Data Output 
ADDRA => ADDRA, -- 14-bit Address Input 
CLKA => CLK, -- Clock 
DIA => ram_3_DIA, -- 4-bit Data Input 
ENA => ENA, -- RAM Enable Input 
WEA => WEA, -- Write Enable Input 
DOB => ram_3_DOB, -- 4-bit Data Output 
ADDRB => ADDRB, -- 12-bit Address Input 
CLKB => CLK, -- Clock 
SSRA => '0', 
SSRB => '0', 
DIB => ram_3_DIB, -- 4-bit Data Input 
ENB => ENB, -- RAM Enable Input 
WEB => WEB -- Write Enable Input 
);
RAM_4_inst : RAMB16_S4_S4 
generic map ( 
INIT_00 => X"0000019b03c2ab170000019b003050d100d000e3000b00130000001800000018",
INIT_01 => X"00030091000180910660010f000c423b00000007000000650000000000000000",
INIT_02 => X"0e2d7405000000100000001000003383000a701300000635000000c300000011",
INIT_03 => X"000000eb00000000000000b8000000000000000900000100000000021c5ae805",
INIT_04 => X"a2828004108581f52aceabc1810820cc6820cc683ed7925acce02affffffffae",
INIT_05 => X"74b16c5c80f4c430a8c932189915c73dfd90ed1a3ea85b2b0ac75f645bc90102",
INIT_06 => X"a7c8926e55800000b0000000000800000047860422d2a065a340c48000c41029",
INIT_07 => X"911a80000100a0011011488d01713032d7558986a5ce2c4e31e7216816f08000",
INIT_08 => X"8746e189110b68c000dd868a2f033e8d61a280caf9f9effb4101d11a010d1409",
INIT_09 => X"0c2fda0740ba28640440004faf0400c0e0011a23b0280280280d140000000c85",
INIT_0A => X"4430220221604605b1156cd001130320ae2260640622f80abcc02c0320037920",
INIT_0B => X"81818196b61ad50327498e8c3f24e430c3d0c30b160b46f9345b03424424c088",
INIT_0C => X"63423907606347041046b6390411120c6308c72044040000000a081101040401",
INIT_0D => X"00000000000000002060088000000007bde0c2c3dddead91a64402c20a912026",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"000000000000000000000000000000000000000000000000000000000f0f8000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map ( 
DOA => ram_4_DOA, -- 4-bit Data Output 
ADDRA => ADDRA, -- 14-bit Address Input 
CLKA => CLK, -- Clock 
DIA => ram_4_DIA, -- 4-bit Data Input 
ENA => ENA, -- RAM Enable Input 
WEA => WEA, -- Write Enable Input 
DOB => ram_4_DOB, -- 4-bit Data Output 
ADDRB => ADDRB, -- 12-bit Address Input 
CLKB => CLK, -- Clock 
SSRA => '0', 
SSRB => '0', 
DIB => ram_4_DIB, -- 4-bit Data Input 
ENB => ENB, -- RAM Enable Input 
WEB => WEB -- Write Enable Input 
);
RAM_5_inst : RAMB16_S4_S4 
generic map ( 
INIT_00 => X"0000003f000223170000003f000050d120d300e3000360130000000000000010",
INIT_01 => X"0000009100000091006a01030000429f000008030000000d0000000000000000",
INIT_02 => X"002d540500000000000000100020030300028013000000350000000300000001",
INIT_03 => X"0000002b000000000000000800000000000000010000002000000002005aa805",
INIT_04 => X"a1028405208541c4e4a89ea180c00002600002600384925a0d002a0000000024",
INIT_05 => X"6e21c87080f4c5142c2832881916623b8d94678aa0a81b2c42d45d641e0d0102",
INIT_06 => X"3e40506ec18000003000000000000800021796209213a0642140c00000c40408",
INIT_07 => X"91c280000100289116818889094120321741010701c7851c7cae0d0807900000",
INIT_08 => X"2205c8c5826c408000b826083902320b098208cb31d1dc0300054098118c1061",
INIT_09 => X"4580182702d82065a098025c0e0d80c0a029502700200200204c1000a6008cb6",
INIT_0A => X"002022d068422422a1c56c804822032d91044065a304e01ae0d06a232003c1a0",
INIT_0B => X"01010190b402d6832c45aa087006e0208280820a180205c834c203984588808b",
INIT_0C => X"43c63a07404205881487243a0431640a4218d440880818026982002000100429",
INIT_0D => X"00000000000000020124808000888087bde0e2c717b8a196064001880aa14006",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"000000000000000000000000000000000000000000000000000000000f0f0000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map ( 
DOA => ram_5_DOA, -- 4-bit Data Output 
ADDRA => ADDRA, -- 14-bit Address Input 
CLKA => CLK, -- Clock 
DIA => ram_5_DIA, -- 4-bit Data Input 
ENA => ENA, -- RAM Enable Input 
WEA => WEA, -- Write Enable Input 
DOB => ram_5_DOB, -- 4-bit Data Output 
ADDRB => ADDRB, -- 12-bit Address Input 
CLKB => CLK, -- Clock 
SSRA => '0', 
SSRB => '0', 
DIB => ram_5_DIB, -- 4-bit Data Input 
ENB => ENB, -- RAM Enable Input 
WEB => WEB -- Write Enable Input 
);
RAM_6_inst : RAMB16_S4_S4 
generic map ( 
INIT_00 => X"0000019b03c022170000019b003050d100d000e3000b00130000000000000000",
INIT_01 => X"00030091000180910660010f000c421b00000003000000650000001000000000",
INIT_02 => X"0e2d7405000000100000001000000303000a001300000635000000c300000011",
INIT_03 => X"000000eb0000000000000088000000000000000900000100000000021c5ae805",
INIT_04 => X"22000000000000f4200e83008040204c60204c603dc69258cc002ac000000012",
INIT_05 => X"56a0e81c8454c032aac9101898035531ec80c9183ca859060a87572017c90800",
INIT_06 => X"8751126455820808b0410101011048202142860800d3a221a144400404c00209",
INIT_07 => X"811a8410100480080051000c01712010d7450102a0c2300e110720e845d08208",
INIT_08 => X"1480e5a9500610c2081d85041d093f0161410441a9e98ffa8201a014010a0808",
INIT_09 => X"0c2fd406809410201400212f0700024221041c13b0900900900a080410084403",
INIT_0A => X"4020000a05414414a1156c9125020100a4a0402016a078007c8000010082f921",
INIT_0B => X"01010086b45ad71107410d003f24a8208320820a0c0880e9305a014200208000",
INIT_0C => X"42c21a03404086080080340a0010840440084740480800210402080101082009",
INIT_0D => X"00000000000000017044808800880087bde02043d51ea082a20400c001a14026",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"000000000000000000000000000000000000000000000000000000000f0f0000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map ( 
DOA => ram_6_DOA, -- 4-bit Data Output 
ADDRA => ADDRA, -- 14-bit Address Input 
CLKA => CLK, -- Clock 
DIA => ram_6_DIA, -- 4-bit Data Input 
ENA => ENA, -- RAM Enable Input 
WEA => WEA, -- Write Enable Input 
DOB => ram_6_DOB, -- 4-bit Data Output 
ADDRB => ADDRB, -- 12-bit Address Input 
CLKB => CLK, -- Clock 
SSRA => '0', 
SSRB => '0', 
DIB => ram_6_DIB, -- 4-bit Data Input 
ENB => ENB, -- RAM Enable Input 
WEB => WEB -- Write Enable Input 
);
RAM_7_inst : RAMB16_S4_S4 
generic map ( 
INIT_00 => X"0000000000100040000000000004000430e0a972000395220000001800000018",
INIT_01 => X"0000410400002104004152000000502800000c24000000000000001800000000",
INIT_02 => X"0020050800000018000000180030058200030522000000000000000800000004",
INIT_03 => X"0000000800000000000000020000000000000002000000610000000200400a08",
INIT_04 => X"61815282b042c2818d503460956a8a918a8a918a810002a0080a4c000000001b",
INIT_05 => X"93308c213e56e2db3311916cdc8a5845088b126d41b3e114b328602264127c81",
INIT_06 => X"545ba37539df7d7d3befafafafbbedf5f5b2b76db1031f22063e46bebee29b31",
INIT_07 => X"8a633efafabed56c8b666452a787b09106198582c58adaf8d6d03683e917df7d",
INIT_08 => X"58c216326db4981f7d421986117c41848661864522022802c30c30660e330c34",
INIT_09 => X"b6d00610c1261822db6df5a05456df1f2fb6a61847d87d87d8330c3edb7d645a",
INIT_0A => X"a6b0916cb66196193060026fb6db0916dadb6122d8db42ad412ab55917dc824f",
INIT_0B => X"8585848803e006f9101a518500310c30c230c30b097cc209bb23096d22d6c245",
INIT_0C => X"60d35b0b6160c0ac2ac2c61b0a9ab615614d68616c2c2df5b6cb7dd9afadf76d",
INIT_0D => X"00000000000000000168008800800807bde0615204502c8b5226aa1aa5b06137",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"000000000000000000000000000000000000000000000000000000000f0f0000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map ( 
DOA => ram_7_DOA, -- 4-bit Data Output 
ADDRA => ADDRA, -- 14-bit Address Input 
CLKA => CLK, -- Clock 
DIA => ram_7_DIA, -- 4-bit Data Input 
ENA => ENA, -- RAM Enable Input 
WEA => WEA, -- Write Enable Input 
DOB => ram_7_DOB, -- 4-bit Data Output 
ADDRB => ADDRB, -- 12-bit Address Input 
CLKB => CLK, -- Clock 
SSRA => '0', 
SSRB => '0', 
DIB => ram_7_DIB, -- 4-bit Data Input 
ENB => ENB, -- RAM Enable Input 
WEB => WEB -- Write Enable Input 
);
end behave;
