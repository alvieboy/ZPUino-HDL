library IEEE;
use IEEE.std_logic_1164.all; 
use IEEE.std_logic_unsigned.all; 
use ieee.numeric_std.all;

entity bootloader_dp_32 is
  port (
    CLK:              in std_logic;
    WEA:  in std_logic;
    ENA:  in std_logic;
    MASKA:    in std_logic_vector(3 downto 0);
    ADDRA:         in std_logic_vector(11 downto 2);
    DIA:        in std_logic_vector(31 downto 0);
    DOA:         out std_logic_vector(31 downto 0);
    WEB:  in std_logic;
    ENB:  in std_logic;
    ADDRB:         in std_logic_vector(11 downto 2);
    DIB:        in std_logic_vector(31 downto 0);
    MASKB:    in std_logic_vector(3 downto 0);
    DOB:         out std_logic_vector(31 downto 0)
  );
end entity bootloader_dp_32;

architecture behave of bootloader_dp_32 is

  subtype RAM_WORD is STD_LOGIC_VECTOR (31 downto 0);
  type RAM_TABLE is array (0 to 1023) of RAM_WORD;
 shared variable RAM: RAM_TABLE := RAM_TABLE'(
x"0b0b0b9b",x"e2040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b9b",x"cc040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fd0608",x"72830609",x"81058205",x"832b2a83",x"ffff0652",x"04000000",x"00000000",x"00000000",x"71fd0608",x"83ffff73",x"83060981",x"05820583",x"2b2b0906",x"7383ffff",x"0b0b0b0b",x"83a70400",x"72098105",x"72057373",x"09060906",x"73097306",x"070a8106",x"53510400",x"00000000",x"00000000",x"72722473",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71737109",x"71068106",x"30720a10",x"0a720a10",x"0a31050a",x"81065151",x"53510400",x"00000000",x"72722673",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"cc040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"720a722b",x"0a535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72729f06",x"0981050b",x"0b0b88af",x"05040000",x"00000000",x"00000000",x"00000000",x"00000000",x"72722aff",x"739f062a",x"0974090a",x"8106ff05",x"06075351",x"04000000",x"00000000",x"00000000",x"71715351",x"020d0406",x"73830609",x"81058205",x"832b0b2b",x"0772fc06",x"0c515104",x"00000000",x"72098105",x"72050970",x"81050906",x"0a810653",x"51040000",x"00000000",x"00000000",x"00000000",x"72098105",x"72050970",x"81050906",x"0a098106",x"53510400",x"00000000",x"00000000",x"00000000",x"71098105",x"52040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72720981",x"05055351",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097206",x"73730906",x"07535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fc0608",x"72830609",x"81058305",x"1010102a",x"81ff0652",x"04000000",x"00000000",x"00000000",x"71fc0608",x"0b0b0b9e",x"ac738306",x"10100508",x"060b0b0b",x"88b20400",x"00000000",x"00000000",x"0b0b0b89",x"80040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"e8040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097081",x"0509060a",x"8106ff05",x"70547106",x"73097274",x"05ff0506",x"07515151",x"04000000",x"72097081",x"0509060a",x"098106ff",x"05705471",x"06730972",x"7405ff05",x"06075151",x"51040000",x"05ff0504",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"810b0b0b",x"0b9f9c0c",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71810552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"02840572",x"10100552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"717105ff",x"05715351",x"020d0400",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"81d53f96",x"853f0400",x"00000000",x"00000000",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101053",x"51047381",x"ff067383",x"06098105",x"83051010",x"102b0772",x"fc060c51",x"51043c04",x"72728072",x"8106ff05",x"09720605",x"71105272",x"0a100a53",x"72ed3851",x"51535104",x"88088c08",x"90087575",x"9d842d50",x"50880856",x"900c8c0c",x"880c5104",x"88088c08",x"90087575",x"9cc92d50",x"50880856",x"900c8c0c",x"880c5104",x"88088c08",x"90088f83",x"2d900c8c",x"0c880c04",x"ff3d0d0b",x"0b0b9fc0",x"3351709e",x"389fa808",x"70085252",x"70802e8a",x"3884129f",x"a80c702d",x"ec39810b",x"0b0b0b9f",x"c034833d",x"0d040480",x"3d0d0b0b",x"0b9ff408",x"802e9738",x"0b0b0b0b",x"800b802e",x"8d380b0b",x"0b9ff451",x"0b0b0bf6",x"873f823d",x"0d0404ff",x"3d0d80c4",x"80808452",x"71087082",x"2a708106",x"51515170",x"f338833d",x"0d04ff3d",x"0d80c480",x"80845271",x"0870812a",x"70810651",x"515170f3",x"38738290",x"0a0c833d",x"0d04fd3d",x"0d755473",x"337081ff",x"06535371",x"802e8e38",x"7281ff06",x"518a9a2d",x"811454e7",x"39853d0d",x"04fe3d0d",x"747080dc",x"8080880c",x"7081ff06",x"ff831154",x"51537181",x"268d3880",x"fd518a9a",x"2d72a032",x"51833972",x"518a9a2d",x"843d0d04",x"fe3d0d74",x"ff175353",x"71ff2e90",x"38727081",x"05543351",x"8add2dff",x"1252ed39",x"843d0d04",x"ff3d0d02",x"8f053352",x"83ffff0b",x"83d00a0c",x"80fe518a",x"9a2d7151",x"8add2d83",x"3d0d04fe",x"3d0d83d0",x"0a087081",x"ff065252",x"8add2d71",x"882a518a",x"dd2d80fe",x"518a9a2d",x"9fd83381",x"05870652",x"719fd834",x"843d0d04",x"fe3d0d9f",x"dc337083",x"2b820781",x"fa065253",x"8bac2d8b",x"cb2d843d",x"0d04fe3d",x"0d9fdc33",x"70832b81",x"0781f906",x"52538bac",x"2d8bcb2d",x"843d0d04",x"82f6ff0b",x"80cc8080",x"880c800b",x"80cc8080",x"840c9f0b",x"83900a0c",x"04ff3d0d",x"73700851",x"5180c880",x"80847008",x"70848080",x"07720c52",x"52833d0d",x"04ff3d0d",x"80c88080",x"84700870",x"fbffff06",x"720c5252",x"833d0d04",x"a0900b80",x"c0800c9f",x"c40b80c0",x"840c9bc3",x"2dff3d0d",x"73518b71",x"0c901152",x"98808072",x"0c80720c",x"700883ff",x"ff06880c",x"833d0d04",x"fa3d0d78",x"7a7dff1e",x"56565855",x"72ff2ea7",x"38805684",x"5275750c",x"74088818",x"0cff1252",x"71f33873",x"84157608",x"720cff15",x"55555272",x"ff2e0981",x"06dd3888",x"3d0d04f9",x"3d0d80d0",x"80808457",x"83d00a0b",x"9ef05258",x"8aba2d8c",x"e12d7651",x"8d892d9f",x"c4708808",x"84299880",x"84057170",x"8405530c",x"5656fb80",x"84a1ad75",x"0c9fac0b",x"88170c80",x"70780c77",x"0c760870",x"83ffff06",x"515683ff",x"ff780ca0",x"80548808",x"53775276",x"518da82d",x"76518cc5",x"2d770855",x"75752e89",x"3880c351",x"8a9a2dff",x"39a08408",x"5574fba0",x"90ae802e",x"893880c2",x"518a9a2d",x"ff399ef8",x"518aba2d",x"80d00a70",x"0870ffbf",x"06720c56",x"5689ff2d",x"8cf82dff",x"3d0d9fd0",x"0881119f",x"d00c5183",x"900a7008",x"70feff06",x"720c5252",x"833d0d04",x"fe3d0d9f",x"d8337083",x"2b818007",x"9fdc3371",x"81f80607",x"5353538b",x"ac2d7481",x"8007518a",x"dd2d8bcb",x"2d843d0d",x"04fe3d0d",x"80d08080",x"84538ce1",x"2d85730c",x"80730c72",x"087081ff",x"06745351",x"528cc52d",x"71880c84",x"3d0d04fc",x"3d0d7653",x"8bf82d81",x"13338214",x"33718180",x"0a297184",x"80802905",x"83163370",x"82802912",x"84183352",x"7105a080",x"05861885",x"19335952",x"53535456",x"54ff1353",x"72ff2e91",x"38737081",x"05553352",x"71757081",x"055734e9",x"3989518f",x"a02d863d",x"0d04f93d",x"0d795680",x"d0808084",x"578ce12d",x"81163382",x"17337182",x"80290553",x"5371802e",x"94388516",x"72555372",x"70810554",x"33770cff",x"145473f3",x"38831633",x"84173371",x"82802905",x"56528054",x"73752797",x"38735877",x"770c7316",x"77085353",x"71733481",x"14547474",x"26ed3876",x"518cc52d",x"9fd83370",x"832b8180",x"079fdc33",x"7181f806",x"07535354",x"8bac2d81",x"84518add",x"2d74882a",x"518add2d",x"74518add",x"2d805473",x"75278f38",x"73167033",x"52528add",x"2d811454",x"ee398bcb",x"2d893d0d",x"04fc3d0d",x"80d08080",x"840b8118",x"54558bf8",x"2d8ce12d",x"86750c74",x"518cc52d",x"8ce12d82",x"750c7270",x"81055433",x"750c7270",x"81055433",x"750c7270",x"81055433",x"750c81ff",x"54727081",x"05543375",x"0cff1454",x"738025f1",x"3874518c",x"c52d8fc9",x"2d880881",x"065271f6",x"38863d0d",x"04fa3d0d",x"785680d0",x"80808454",x"8ce12d86",x"740c7351",x"8cc52d8c",x"e12d81ad",x"740c8116",x"33821733",x"71828029",x"05831833",x"760c8418",x"33760c85",x"1833760c",x"58528055",x"747727af",x"3874802e",x"88388ce1",x"2d81ad74",x"0c741686",x"1133750c",x"87113375",x"0c527351",x"8cc52d8f",x"c92d8808",x"81065271",x"f6388215",x"55ce398c",x"e12d8474",x"0c73518c",x"c52d9fd8",x"3370832b",x"8180079f",x"dc337181",x"f8060753",x"53538bac",x"2d818751",x"8add2d8b",x"cb2d883d",x"0d04fc3d",x"0d768111",x"33821233",x"71902b71",x"882b0783",x"14337072",x"07882b84",x"16337107",x"51525356",x"57555288",x"518fa02d",x"81ff518a",x"9a2d80c4",x"80808454",x"73087081",x"2a708106",x"51515271",x"f3387284",x"80800780",x"c4808084",x"0c863d0d",x"04fd3d0d",x"8fc92d88",x"08880881",x"06535371",x"f3389fd8",x"3370832b",x"8180079f",x"dc337181",x"f8060753",x"53548bac",x"2d818351",x"8add2d72",x"518add2d",x"8bcb2d85",x"3d0d04fb",x"3d0d800b",x"9fd00c80",x"709ebc58",x"55557570",x"84055708",x"5372802e",x"8a388114",x"81712b76",x"07565381",x"14548c74",x"27e4389f",x"d8337083",x"2b818007",x"9fdc3371",x"81f80607",x"5354548b",x"ac2d8181",x"518add2d",x"94529fac",x"518b8c2d",x"94529fac",x"518b8c2d",x"74982a51",x"8add2d74",x"902a518a",x"dd2d7488",x"2a518add",x"2d74518a",x"dd2d8bcb",x"2d873d0d",x"04fe3d0d",x"800b9fd0",x"0c9fd833",x"70832b81",x"80079fdc",x"337181f8",x"06075353",x"538bac2d",x"8182518a",x"dd2d80d0",x"80808452",x"8ce12d81",x"f90a0b80",x"d080809c",x"0c710872",x"52538cc5",x"2d729fe0",x"0c72902a",x"518add2d",x"9fe00888",x"2a518add",x"2d9fe008",x"518add2d",x"8fc92d88",x"08518add",x"2d8bcb2d",x"843d0d04",x"803d0d81",x"0b9fd40c",x"800b8390",x"0a0c8551",x"8fa02d82",x"3d0d0480",x"3d0d800b",x"9fd40c8c",x"ac2d8651",x"8fa02d82",x"3d0d04fd",x"3d0d80d0",x"80808454",x"8a518fa0",x"2d8ce12d",x"9fc47452",x"538d892d",x"72880884",x"29988084",x"05717084",x"05530c52",x"fb8084a1",x"ad720c9f",x"ac0b8814",x"0c73518c",x"c52d89ff",x"2d8cf82d",x"ffb23d0d",x"80d23d08",x"56800b9f",x"d40c800b",x"9fd00c80",x"0bdf8017",x"9fb17190",x"2a715656",x"57555772",x"72708105",x"54347388",x"2a537272",x"34738216",x"3475982a",x"52718b16",x"3475902a",x"52718c16",x"3475882a",x"52718d16",x"34758e16",x"348f830b",x"80c0800c",x"8480b30b",x"80c48080",x"840c80c8",x"8080a453",x"fbffff73",x"08707206",x"750c5354",x"80c88080",x"94700870",x"7606720c",x"5353880b",x"80c08080",x"840c810b",x"900a0c9f",x"90518aba",x"2d8cac2d",x"fe88880b",x"80dc8080",x"840c81f2",x"0b80d00a",x"0c80d080",x"80847052",x"528cc52d",x"8ce12d71",x"518cc52d",x"8ce12d84",x"720c7151",x"8cc52d76",x"77565480",x"c4808084",x"08708106",x"5152719e",x"389fd408",x"5372ec38",x"9fd00852",x"87e87227",x"e2387290",x"0a0c7283",x"900a0c9b",x"bb2d8290",x"0a085374",x"802e81c9",x"387280fe",x"2e098106",x"81823876",x"802effbb",x"38805582",x"7727ffb3",x"3883d00a",x"08527175",x"2e098106",x"b738883d",x"3370872a",x"81325353",x"71802e97",x"38728706",x"5271ff8f",x"38749fdc",x"34749fd8",x"348bf82d",x"ff813972",x"b8067083",x"2a9fdc33",x"55515271",x"732e8738",x"8c922dfe",x"ea398113",x"87065271",x"9fdc3402",x"9d053352",x"718d26fe",x"d6387184",x"299eb805",x"80d13dfd",x"e1055270",x"08515271",x"2dfec039",x"7280fd2e",x"09810686",x"388154fe",x"b2397682",x"9f26a538",x"73802e87",x"388073a0",x"32545472",x"80dc8080",x"880c80d0",x"3d7705fd",x"e0055272",x"72348117",x"57fe8839",x"8055fe83",x"397280fe",x"2e098106",x"fdf93874",x"57ff0b83",x"d00a0c81",x"775555fd",x"ea39ff3d",x"0d9c9d2d",x"73528051",x"97c82d83",x"3d0d0483",x"fffff80d",x"8de30483",x"fffff80d",x"80c08804",x"880880c0",x"80808808",x"80c08008",x"2d50880c",x"810b900a",x"0c048070",x"0cfaad95",x"b4da0b81",x"80807171",x"0c718008",x"2e873870",x"11519bee",x"04519baa",x"2d000000",x"00000000",x"00000000",x"00000000",x"820b80c0",x"8080900c",x"0b0b0b04",x"0083f00a",x"0b800ba0",x"80721208",x"720c8412",x"5271712e",x"ff05f238",x"028c050d",x"9c900400",x"00000000",x"00000000",x"00000000",x"00fb3d0d",x"77795555",x"80567476",x"25863874",x"30558156",x"73802588",x"38733076",x"81325754",x"80537352",x"745180ca",x"3f880854",x"75802e85",x"38880830",x"5473880c",x"873d0d04",x"fa3d0d78",x"7a575580",x"57747725",x"86387430",x"55815775",x"9f2c5481",x"53757432",x"74315274",x"51943f88",x"08547680",x"2e853888",x"08305473",x"880c883d",x"0d04fc3d",x"0d767853",x"54815380",x"55873971",x"10731054",x"52737226",x"5172802e",x"a7387080",x"2e863871",x"8025e838",x"72802e98",x"38717426",x"89387372",x"31757407",x"56547281",x"2a72812a",x"5353e539",x"73517883",x"38745170",x"880c863d",x"0d04ff3d",x"0d9fe80b",x"fc055271",x"08ff2e8b",x"38710851",x"702dfc12",x"52f13983",x"3d0d0404",x"eafe3f04",x"00ffffff",x"ff00ffff",x"ffff00ff",x"ffffff00",x"00000a77",x"00000af1",x"00000a3d",x"00000846",x"00000b5c",x"00000b73",x"0000094d",x"000009ea",x"000007ef",x"00000b87",x"000008ed",x"00000000",x"00000000",x"43500d0a",x"00000000",x"4c6f6164",x"65642c20",x"73746172",x"74696e67",x"2e2e2e0d",x"0a000000",x"0d0a5a50",x"55494e4f",x"0d0a0000",x"00000000",x"00000000",x"00000000",x"00000ff0",x"02010600",x"00000000",x"05b8d800",x"b4041700",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"ffffffff",x"00000000",x"ffffffff",x"00000000",x"00000000",x"00000000",x"00000000");

begin

  process (clk)
  begin
    if rising_edge(clk) then
      if ENA='1' then
        if WEA='1' then
          RAM(conv_integer(ADDRA) ) := DIA;
        end if;
        DOA <= RAM(conv_integer(ADDRA)) ;
      end if;
    end if;
  end process;  

  process (clk)
  begin
    if rising_edge(clk) then
      if ENB='1' then
        if WEB='1' then
          RAM( conv_integer(ADDRB) ) := DIB;
        end if;
        DOB <= RAM(conv_integer(ADDRB)) ;
      end if;
    end if;
  end process;  
end behave;
