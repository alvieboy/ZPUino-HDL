library IEEE;
use IEEE.std_logic_1164.all; 
use IEEE.std_logic_unsigned.all; 
use ieee.numeric_std.all;

entity bootloader_dp_32 is
  port (
    CLK:              in std_logic;
    WEA:  in std_logic;
    ENA:  in std_logic;
    MASKA:    in std_logic_vector(3 downto 0);
    ADDRA:         in std_logic_vector(11 downto 2);
    DIA:        in std_logic_vector(31 downto 0);
    DOA:         out std_logic_vector(31 downto 0);
    WEB:  in std_logic;
    ENB:  in std_logic;
    ADDRB:         in std_logic_vector(11 downto 2);
    DIB:        in std_logic_vector(31 downto 0);
    MASKB:    in std_logic_vector(3 downto 0);
    DOB:         out std_logic_vector(31 downto 0)
  );
end entity bootloader_dp_32;

architecture behave of bootloader_dp_32 is

  subtype RAM_WORD is STD_LOGIC_VECTOR (31 downto 0);
  type RAM_TABLE is array (0 to 1023) of RAM_WORD;
 shared variable RAM: RAM_TABLE := RAM_TABLE'(
x"0b0b0b98",x"96040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b98",x"b2040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fd0608",x"72830609",x"81058205",x"832b2a83",x"ffff0652",x"04000000",x"00000000",x"00000000",x"71fd0608",x"83ffff73",x"83060981",x"05820583",x"2b2b0906",x"7383ffff",x"0b0b0b0b",x"83a70400",x"72098105",x"72057373",x"09060906",x"73097306",x"070a8106",x"53510400",x"00000000",x"00000000",x"72722473",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71737109",x"71068106",x"30720a10",x"0a720a10",x"0a31050a",x"81065151",x"53510400",x"00000000",x"72722673",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"c3040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"720a722b",x"0a535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72729f06",x"0981050b",x"0b0b88a6",x"05040000",x"00000000",x"00000000",x"00000000",x"00000000",x"72722aff",x"739f062a",x"0974090a",x"8106ff05",x"06075351",x"04000000",x"00000000",x"00000000",x"71715351",x"020d0406",x"73830609",x"81058205",x"832b0b2b",x"0772fc06",x"0c515104",x"00000000",x"72098105",x"72050970",x"81050906",x"0a810653",x"51040000",x"00000000",x"00000000",x"00000000",x"72098105",x"72050970",x"81050906",x"0a098106",x"53510400",x"00000000",x"00000000",x"00000000",x"71098105",x"52040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72720981",x"05055351",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097206",x"73730906",x"07535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fc0608",x"72830609",x"81058305",x"1010102a",x"81ff0652",x"04000000",x"00000000",x"00000000",x"71fc0608",x"0b0b0b9e",x"88738306",x"10100508",x"060b0b0b",x"88a90400",x"00000000",x"00000000",x"0b0b0b88",x"f7040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"df040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097081",x"0509060a",x"8106ff05",x"70547106",x"73097274",x"05ff0506",x"07515151",x"04000000",x"72097081",x"0509060a",x"098106ff",x"05705471",x"06730972",x"7405ff05",x"06075151",x"51040000",x"05ff0504",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"810b0b0b",x"0b9ed00c",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71810552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"02840572",x"10100552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"717105ff",x"05715351",x"020d0400",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"81d43f95",x"d83f0410",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10105351",x"047381ff",x"06738306",x"09810583",x"05101010",x"2b0772fc",x"060c5151",x"043c0472",x"72807281",x"06ff0509",x"72060571",x"1052720a",x"100a5372",x"ed385151",x"53510488",x"088c0890",x"08757599",x"8b2d5050",x"88085690",x"0c8c0c88",x"0c510488",x"088c0890",x"08757598",x"c72d5050",x"88085690",x"0c8c0c88",x"0c510488",x"088c0890",x"088df62d",x"900c8c0c",x"880c04ff",x"3d0d0b0b",x"0b9ee033",x"5170a638",x"9edc0870",x"08525270",x"802e9238",x"84129edc",x"0c702d9e",x"dc087008",x"525270f0",x"38810b0b",x"0b0b9ee0",x"34833d0d",x"0404803d",x"0d0b0b0b",x"9f8c0880",x"2e8e380b",x"0b0b0b80",x"0b802e09",x"81068538",x"823d0d04",x"0b0b0b9f",x"8c510b0b",x"0bf6813f",x"823d0d04",x"04ff3d0d",x"80c48080",x"84527108",x"70822a70",x"81065151",x"5170f338",x"833d0d04",x"ff3d0d80",x"c4808084",x"52710870",x"812a7081",x"06515151",x"70f33873",x"82900a0c",x"833d0d04",x"fe3d0d74",x"7080dc80",x"80880c70",x"81ff06ff",x"83115451",x"53718126",x"8d3880fd",x"518aa02d",x"72a03251",x"83397251",x"8aa02d84",x"3d0d0480",x"3d0d83ff",x"ff0b83d0",x"0a0c80fe",x"518aa02d",x"823d0d04",x"ff3d0d83",x"d00a0870",x"882a5252",x"8ac02d71",x"81ff0651",x"8ac02d80",x"fe518aa0",x"2d833d0d",x"0482f6ff",x"0b80cc80",x"80880c80",x"0b80cc80",x"80840c9f",x"0b83900a",x"0c04ff3d",x"0d737008",x"515180c8",x"80808470",x"08708480",x"8007720c",x"5252833d",x"0d04ff3d",x"0d80c880",x"80847008",x"70fbffff",x"06720c52",x"52833d0d",x"04a0900b",x"a0800c9e",x"e40ba084",x"0c98ab2d",x"ff3d0d73",x"518b710c",x"90115291",x"c080720c",x"80720c70",x"0883ffff",x"06880c83",x"3d0d04fa",x"3d0d787a",x"7dff1e57",x"57585373",x"ff2ea738",x"80568452",x"75730c72",x"0888180c",x"ff125271",x"f3387484",x"16740872",x"0cff1656",x"565273ff",x"2e098106",x"dd38883d",x"0d04f83d",x"0d80d080",x"80845783",x"d00a598b",x"da2d7651",x"8c802d9e",x"e4708808",x"101091c0",x"84057170",x"8405530c",x"5656fb80",x"84a1ad75",x"0c9ec00b",x"88170c80",x"70780c77",x"0c760883",x"ffff0656",x"81df800b",x"88082783",x"38ff3983",x"ffff790c",x"a0805488",x"08537852",x"76518c9f",x"2d76518b",x"be2d7808",x"5574762e",x"893880c3",x"518aa02d",x"ff39a084",x"085574fb",x"a0849e80",x"2e893880",x"c2518aa0",x"2dff3980",x"d00a7008",x"70ffbf06",x"720c5656",x"8a852d8b",x"f12dff3d",x"0d9ef008",x"81119ef0",x"0c518390",x"0a700870",x"feff0672",x"0c525283",x"3d0d0480",x"3d0d8aef",x"2d728180",x"07518ac0",x"2d8b842d",x"823d0d04",x"fe3d0d80",x"d0808084",x"538bda2d",x"85730c80",x"730c7208",x"7081ff06",x"74535152",x"8bbe2d71",x"880c843d",x"0d04fc3d",x"0d768111",x"33821233",x"7181800a",x"29718480",x"80290583",x"14337082",x"80291284",x"16335271",x"05a08005",x"86168517",x"33575253",x"53555755",x"53ff1353",x"72ff2e91",x"38737081",x"05553352",x"71757081",x"055734e9",x"3989518e",x"932d863d",x"0d04f93d",x"0d795780",x"d0808084",x"568bda2d",x"81173382",x"18337182",x"80290553",x"5371802e",x"94388517",x"72555372",x"70810554",x"33760cff",x"145473f3",x"38831733",x"84183371",x"82802905",x"56528054",x"73752797",x"38735877",x"760c7317",x"76085353",x"71733481",x"14547474",x"26ed3875",x"518bbe2d",x"8aef2d81",x"84518ac0",x"2d74882a",x"518ac02d",x"74518ac0",x"2d805473",x"75278f38",x"73177033",x"52528ac0",x"2d811454",x"ee398b84",x"2d893d0d",x"04f93d0d",x"795680d0",x"80808455",x"8bda2d86",x"750c7451",x"8bbe2d8b",x"da2d81ad",x"70760c81",x"17338218",x"33718280",x"29058319",x"33780c84",x"1933780c",x"85193378",x"0c595353",x"80547377",x"27b33872",x"5873802e",x"87388bda",x"2d77750c",x"73168611",x"33760c87",x"1133760c",x"5274518b",x"be2d8ea8",x"2d880881",x"065271f6",x"38821454",x"767426d1",x"388bda2d",x"84750c74",x"518bbe2d",x"8aef2d81",x"87518ac0",x"2d8b842d",x"893d0d04",x"fc3d0d76",x"81113382",x"12337190",x"2b71882b",x"07831433",x"70720788",x"2b841633",x"71075152",x"53575754",x"5288518e",x"932d81ff",x"518aa02d",x"80c48080",x"84537208",x"70812a70",x"81065151",x"5271f338",x"73848080",x"0780c480",x"80840c86",x"3d0d04fe",x"3d0d8ea8",x"2d880888",x"08810653",x"5371f338",x"8aef2d81",x"83518ac0",x"2d72518a",x"c02d8b84",x"2d843d0d",x"04fe3d0d",x"800b9ef0",x"0c8aef2d",x"8181518a",x"c02d9ec0",x"538f5272",x"70810554",x"33518ac0",x"2dff1252",x"71ff2e09",x"8106ec38",x"8b842d84",x"3d0d04fe",x"3d0d800b",x"9ef00c8a",x"ef2d8182",x"518ac02d",x"80d08080",x"84528bda",x"2d81f90a",x"0b80d080",x"809c0c71",x"08725253",x"8bbe2d72",x"9ef80c72",x"902a518a",x"c02d9ef8",x"08882a51",x"8ac02d9e",x"f808518a",x"c02d8ea8",x"2d880851",x"8ac02d8b",x"842d843d",x"0d04803d",x"0d810b9e",x"f40c800b",x"83900a0c",x"85518e93",x"2d823d0d",x"04803d0d",x"800b9ef4",x"0c8ba52d",x"86518e93",x"2d823d0d",x"04fd3d0d",x"80d08080",x"84548a51",x"8e932d8b",x"da2d9ee4",x"7452538c",x"802d7288",x"08101091",x"c0840571",x"70840553",x"0c52fb80",x"84a1ad72",x"0c9ec00b",x"88140c73",x"518bbe2d",x"8a852d8b",x"f12dfc3d",x"0d80d080",x"80847052",x"558bbe2d",x"8bda2d8b",x"750c7680",x"d0808094",x"0c80750c",x"a0805477",x"5383d00a",x"5274518c",x"9f2d7451",x"8bbe2d8a",x"852d8bf1",x"2dffab3d",x"0d800b9e",x"f40c800b",x"9ef00c80",x"0b8df60b",x"a0800c57",x"80c48080",x"84558480",x"b3750c80",x"c88080a4",x"53fbffff",x"73087072",x"06750c53",x"5480c880",x"80947008",x"70760672",x"0c5353a8",x"7099c371",x"70840553",x"0c9aa071",x"0c539bb9",x"0b88120c",x"9cc80b8c",x"120c94b2",x"0b90120c",x"53880b80",x"c0808084",x"0c900a53",x"81730c8b",x"a52dfe88",x"880b80dc",x"8080840c",x"81f20b80",x"d00a0c80",x"d0808084",x"7052528b",x"be2d8bda",x"2d71518b",x"be2d8bda",x"2d84720c",x"71518bbe",x"2d767776",x"75933d41",x"415b5b5b",x"83d00a5c",x"78087081",x"06515271",x"9d389ef4",x"085372f0",x"389ef008",x"5287e872",x"27e63872",x"7e0c7283",x"900a0c98",x"a42d8290",x"0a085379",x"802e81b4",x"387280fe",x"2e098106",x"80f43876",x"802ec138",x"807d7858",x"565a8277",x"27ffb538",x"83ffff7c",x"0c79fe18",x"53537972",x"27983880",x"dc808088",x"72555872",x"15703379",x"0c528113",x"53737326",x"f238ff16",x"75115475",x"05ff0570",x"33743370",x"72882b07",x"7f085351",x"55515271",x"732e0981",x"06feed38",x"74335372",x"8a26fee4",x"38721010",x"9e940575",x"52700851",x"52712dfe",x"d3397280",x"fd2e0981",x"06863881",x"5bfec539",x"76829f26",x"9e387a80",x"2e873880",x"73a03254",x"5b80d73d",x"7705fde0",x"05527272",x"34811757",x"fea23980",x"5afe9d39",x"7280fe2e",x"098106fe",x"93387957",x"ff7c0c81",x"775c5afe",x"8739ff3d",x"0d805280",x"5194e92d",x"833d0d04",x"81fff80d",x"8cda0481",x"fff80da0",x"88048808",x"80c08080",x"8808a080",x"082d5088",x"0c810b90",x"0a0c04fb",x"3d0d7779",x"55558056",x"757524ab",x"38807424",x"9d388053",x"73527451",x"80e13f88",x"08547580",x"2e853888",x"08305473",x"880c873d",x"0d047330",x"76813257",x"54dc3974",x"30558156",x"738025d2",x"38ec39fa",x"3d0d787a",x"57558057",x"767524a4",x"38759f2c",x"54815375",x"74327431",x"5274519b",x"3f880854",x"76802e85",x"38880830",x"5473880c",x"883d0d04",x"74305581",x"57d739fc",x"3d0d7678",x"53548153",x"80747326",x"52557280",x"2e983870",x"802ea938",x"807224a4",x"38711073",x"10757226",x"53545272",x"ea387351",x"78833874",x"5170880c",x"863d0d04",x"72812a72",x"812a5353",x"72802ee6",x"38717426",x"ef387372",x"31757407",x"74812a74",x"812a5555",x"5654e539",x"fc3d0d76",x"70797b55",x"5555558f",x"72278c38",x"72750783",x"06517080",x"2ea738ff",x"125271ff",x"2e983872",x"70810554",x"33747081",x"055634ff",x"125271ff",x"2e098106",x"ea387488",x"0c863d0d",x"04745172",x"70840554",x"08717084",x"05530c72",x"70840554",x"08717084",x"05530c72",x"70840554",x"08717084",x"05530c72",x"70840554",x"08717084",x"05530cf0",x"1252718f",x"26c93883",x"72279538",x"72708405",x"54087170",x"8405530c",x"fc125271",x"8326ed38",x"7054ff83",x"39fc3d0d",x"76797102",x"8c059f05",x"33575553",x"55837227",x"8a387483",x"06517080",x"2ea238ff",x"125271ff",x"2e933873",x"73708105",x"5534ff12",x"5271ff2e",x"098106ef",x"3874880c",x"863d0d04",x"7474882b",x"75077071",x"902b0751",x"54518f72",x"27a53872",x"71708405",x"530c7271",x"70840553",x"0c727170",x"8405530c",x"72717084",x"05530cf0",x"1252718f",x"26dd3883",x"72279038",x"72717084",x"05530cfc",x"12527183",x"26f23870",x"53ff9039",x"fb3d0d77",x"79707207",x"83065354",x"52709338",x"71737308",x"54565471",x"73082e80",x"c4387375",x"54527133",x"7081ff06",x"52547080",x"2e9d3872",x"33557075",x"2e098106",x"95388112",x"81147133",x"7081ff06",x"54565452",x"70e53872",x"33557381",x"ff067581",x"ff067171",x"31880c52",x"52873d0d",x"04710970",x"f7fbfdff",x"140670f8",x"84828180",x"06515151",x"70973884",x"14841671",x"08545654",x"7175082e",x"dc387375",x"5452ff96",x"39800b88",x"0c873d0d",x"04ff3d0d",x"9f800bfc",x"05700852",x"5270ff2e",x"9138702d",x"fc127008",x"525270ff",x"2e098106",x"f138833d",x"0d0404eb",x"9a3f0400",x"00ffffff",x"ff00ffff",x"ffff00ff",x"ffffff00",x"0000093d",x"0000096f",x"00000917",x"000007a2",x"000009c6",x"000009dd",x"00000835",x"000008c4",x"0000074e",x"000009f1",x"01090460",x"00006f80",x"05b8d800",x"b4010f00",x"00000000",x"00000000",x"00000000",x"00000f88",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"ffffffff",x"00000000",x"ffffffff",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000");

begin

  process (clk)
  begin
    if rising_edge(clk) then
      if ENA='1' then
        if WEA='1' then
          RAM(conv_integer(ADDRA) ) := DIA;
        end if;
        DOA <= RAM(conv_integer(ADDRA)) ;
      end if;
    end if;
  end process;  

  process (clk)
  begin
    if rising_edge(clk) then
      if ENB='1' then
        if WEB='1' then
          RAM( conv_integer(ADDRB) ) := DIB;
        end if;
        DOB <= RAM(conv_integer(ADDRB)) ;
      end if;
    end if;
  end process;  
end behave;
