library IEEE;
use IEEE.std_logic_1164.all; 
use IEEE.std_logic_unsigned.all; 
use ieee.numeric_std.all;

entity bootloader_dp_32 is
  port (
    CLK:              in std_logic;
    WEA:  in std_logic;
    ENA:  in std_logic;
    MASKA:    in std_logic_vector(3 downto 0);
    ADDRA:         in std_logic_vector(11 downto 2);
    DIA:        in std_logic_vector(31 downto 0);
    DOA:         out std_logic_vector(31 downto 0);
    WEB:  in std_logic;
    ENB:  in std_logic;
    ADDRB:         in std_logic_vector(11 downto 2);
    DIB:        in std_logic_vector(31 downto 0);
    MASKB:    in std_logic_vector(3 downto 0);
    DOB:         out std_logic_vector(31 downto 0)
  );
end entity bootloader_dp_32;

architecture behave of bootloader_dp_32 is

  subtype RAM_WORD is STD_LOGIC_VECTOR (31 downto 0);
  type RAM_TABLE is array (0 to 1023) of RAM_WORD;
 shared variable RAM: RAM_TABLE := RAM_TABLE'(
x"0b0b0b98",x"c3040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b98",x"ae040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fd0608",x"72830609",x"81058205",x"832b2a83",x"ffff0652",x"04000000",x"00000000",x"00000000",x"71fd0608",x"83ffff73",x"83060981",x"05820583",x"2b2b0906",x"7383ffff",x"0b0b0b0b",x"83a70400",x"72098105",x"72057373",x"09060906",x"73097306",x"070a8106",x"53510400",x"00000000",x"00000000",x"72722473",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71737109",x"71068106",x"30720a10",x"0a720a10",x"0a31050a",x"81065151",x"53510400",x"00000000",x"72722673",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"c3040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"720a722b",x"0a535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72729f06",x"0981050b",x"0b0b88a6",x"05040000",x"00000000",x"00000000",x"00000000",x"00000000",x"72722aff",x"739f062a",x"0974090a",x"8106ff05",x"06075351",x"04000000",x"00000000",x"00000000",x"71715351",x"020d0406",x"73830609",x"81058205",x"832b0b2b",x"0772fc06",x"0c515104",x"00000000",x"72098105",x"72050970",x"81050906",x"0a810653",x"51040000",x"00000000",x"00000000",x"00000000",x"72098105",x"72050970",x"81050906",x"0a098106",x"53510400",x"00000000",x"00000000",x"00000000",x"71098105",x"52040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72720981",x"05055351",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097206",x"73730906",x"07535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fc0608",x"72830609",x"81058305",x"1010102a",x"81ff0652",x"04000000",x"00000000",x"00000000",x"71fc0608",x"0b0b0b9a",x"e8738306",x"10100508",x"060b0b0b",x"88a90400",x"00000000",x"00000000",x"0b0b0b88",x"f7040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"df040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097081",x"0509060a",x"8106ff05",x"70547106",x"73097274",x"05ff0506",x"07515151",x"04000000",x"72097081",x"0509060a",x"098106ff",x"05705471",x"06730972",x"7405ff05",x"06075151",x"51040000",x"05ff0504",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"810b0b0b",x"0b9bcc0c",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71810552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"02840572",x"10100552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"717105ff",x"05715351",x"020d0400",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"81d43f92",x"b63f0410",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10105351",x"047381ff",x"06738306",x"09810583",x"05101010",x"2b0772fc",x"060c5151",x"043c0472",x"72807281",x"06ff0509",x"72060571",x"1052720a",x"100a5372",x"ed385151",x"53510488",x"088c0890",x"08757599",x"a62d5050",x"88085690",x"0c8c0c88",x"0c510488",x"088c0890",x"08757598",x"e22d5050",x"88085690",x"0c8c0c88",x"0c510488",x"088c0890",x"088e9d2d",x"900c8c0c",x"880c04ff",x"3d0d0b0b",x"0b9bf033",x"5170a638",x"9bd80870",x"08525270",x"802e9238",x"84129bd8",x"0c702d9b",x"d8087008",x"525270f0",x"38810b0b",x"0b0b9bf0",x"34833d0d",x"0404803d",x"0d0b0b0b",x"9c9c0880",x"2e8e380b",x"0b0b0b80",x"0b802e09",x"81068538",x"823d0d04",x"0b0b0b9c",x"9c510b0b",x"0bf6813f",x"823d0d04",x"04ff3d0d",x"80c48080",x"84527108",x"70822a70",x"81065151",x"5170f338",x"833d0d04",x"ff3d0d80",x"c4808084",x"52710870",x"812a7081",x"06515151",x"70f33873",x"82900a0c",x"833d0d04",x"fd3d0d75",x"54733370",x"81ff0653",x"5371802e",x"8e387281",x"ff06518a",x"a02d8114",x"54e73985",x"3d0d04fe",x"3d0d7470",x"80dc8080",x"880c7081",x"ff06ff83",x"11545153",x"7181268d",x"3880fd51",x"8aa02d72",x"a0325183",x"3972518a",x"a02d843d",x"0d04803d",x"0d83ffff",x"0b83d00a",x"0c80fe51",x"8aa02d82",x"3d0d04ff",x"3d0d83d0",x"0a087088",x"2a52528a",x"e32d7181",x"ff06518a",x"e32d80fe",x"518aa02d",x"833d0d04",x"82f6ff0b",x"80cc8080",x"880c800b",x"80cc8080",x"840c9f0b",x"83900a0c",x"04ff3d0d",x"73700851",x"5180c880",x"80847008",x"70848080",x"07720c52",x"52833d0d",x"04ff3d0d",x"80c88080",x"84700870",x"fbffff06",x"720c5252",x"833d0d04",x"a0900ba0",x"800c9bf4",x"0ba0840c",x"98a72dff",x"3d0d7351",x"8b710c90",x"115291c0",x"80720c80",x"720c7008",x"83ffff06",x"880c833d",x"0d04fa3d",x"0d787a7d",x"ff1e5757",x"585373ff",x"2ea73880",x"56845275",x"730c7208",x"88180cff",x"125271f3",x"38748416",x"7408720c",x"ff165656",x"5273ff2e",x"098106dd",x"38883d0d",x"04f93d0d",x"80d08080",x"845683d0",x"0a0b9ba0",x"52588ac0",x"2d8bfd2d",x"75518ca3",x"2d9bf470",x"88081010",x"91c08405",x"71708405",x"530c5657",x"fb8084a1",x"ad750c9b",x"dc0b8818",x"0c807077",x"0c760c75",x"087083ff",x"ff065157",x"83ffff78",x"0ca08054",x"88085377",x"5275518c",x"c22d7551",x"8be12d77",x"08557477",x"2e893880",x"c3518aa0",x"2dff39a0",x"84085574",x"fba0849e",x"802e8938",x"80c2518a",x"a02dff39",x"9ba8518a",x"c02d80d0",x"0a700870",x"ffbf0672",x"0c56568a",x"852d8c94",x"2dff3d0d",x"9c800881",x"119c800c",x"5183900a",x"700870fe",x"ff06720c",x"5252833d",x"0d04803d",x"0d8b922d",x"72818007",x"518ae32d",x"8ba72d82",x"3d0d04fe",x"3d0d80d0",x"80808453",x"8bfd2d85",x"730c8073",x"0c720870",x"81ff0674",x"5351528b",x"e12d7188",x"0c843d0d",x"04fc3d0d",x"76811133",x"82123371",x"81800a29",x"71848080",x"29058314",x"33708280",x"29128416",x"33527105",x"a0800586",x"16851733",x"57525353",x"55575553",x"ff135372",x"ff2e9138",x"73708105",x"55335271",x"75708105",x"5734e939",x"89518eba",x"2d863d0d",x"04f93d0d",x"795780d0",x"80808456",x"8bfd2d81",x"17338218",x"33718280",x"29055353",x"71802e94",x"38851772",x"55537270",x"81055433",x"760cff14",x"5473f338",x"83173384",x"18337182",x"80290556",x"52805473",x"75279738",x"73587776",x"0c731776",x"08535371",x"73348114",x"54747426",x"ed387551",x"8be12d8b",x"922d8184",x"518ae32d",x"74882a51",x"8ae32d74",x"518ae32d",x"80547375",x"278f3873",x"17703352",x"528ae32d",x"811454ee",x"398ba72d",x"893d0d04",x"f93d0d79",x"5680d080",x"8084558b",x"fd2d8675",x"0c74518b",x"e12d8bfd",x"2d81ad70",x"760c8117",x"33821833",x"71828029",x"05831933",x"780c8419",x"33780c85",x"1933780c",x"59535380",x"54737727",x"b3387258",x"73802e87",x"388bfd2d",x"77750c73",x"16861133",x"760c8711",x"33760c52",x"74518be1",x"2d8ecf2d",x"88088106",x"5271f638",x"82145476",x"7426d138",x"8bfd2d84",x"750c7451",x"8be12d8b",x"922d8187",x"518ae32d",x"8ba72d89",x"3d0d04fc",x"3d0d7681",x"11338212",x"3371902b",x"71882b07",x"83143370",x"7207882b",x"84163371",x"07515253",x"57575452",x"88518eba",x"2d81ff51",x"8aa02d80",x"c4808084",x"53720870",x"812a7081",x"06515152",x"71f33873",x"84808007",x"80c48080",x"840c863d",x"0d04fe3d",x"0d8ecf2d",x"88088808",x"81065353",x"71f3388b",x"922d8183",x"518ae32d",x"72518ae3",x"2d8ba72d",x"843d0d04",x"fe3d0d80",x"0b9c800c",x"8b922d81",x"81518ae3",x"2d9bdc53",x"93527270",x"81055433",x"518ae32d",x"ff125271",x"ff2e0981",x"06ec388b",x"a72d843d",x"0d04fe3d",x"0d800b9c",x"800c8b92",x"2d818251",x"8ae32d80",x"d0808084",x"528bfd2d",x"81f90a0b",x"80d08080",x"9c0c7108",x"7252538b",x"e12d729c",x"880c7290",x"2a518ae3",x"2d9c8808",x"882a518a",x"e32d9c88",x"08518ae3",x"2d8ecf2d",x"8808518a",x"e32d8ba7",x"2d843d0d",x"04803d0d",x"810b9c84",x"0c800b83",x"900a0c85",x"518eba2d",x"823d0d04",x"803d0d80",x"0b9c840c",x"8bc82d86",x"518eba2d",x"823d0d04",x"fd3d0d80",x"d0808084",x"548a518e",x"ba2d8bfd",x"2d9bf474",x"52538ca3",x"2d728808",x"101091c0",x"84057170",x"8405530c",x"52fb8084",x"a1ad720c",x"9bdc0b88",x"140c7351",x"8be12d8a",x"852d8c94",x"2dffab3d",x"0d80d93d",x"0856800b",x"9c840c80",x"0b9c800c",x"800bdf80",x"179be171",x"902a7156",x"56575557",x"72727081",x"05543473",x"882a5372",x"72347382",x"1634758b",x"16348e9d",x"0ba0800c",x"80c48080",x"84558480",x"b3750c80",x"c88080a4",x"53fbffff",x"73087072",x"06750c53",x"5480c880",x"80947008",x"70760672",x"0c535388",x"0b80c080",x"80840c90",x"0a538173",x"0c9bc051",x"8ac02d8b",x"c82dfe88",x"880b80dc",x"8080840c",x"81f20b80",x"d00a0c80",x"d0808084",x"7052528b",x"e12d8bfd",x"2d71518b",x"e12d8bfd",x"2d84720c",x"71518be1",x"2d767776",x"75933d41",x"415b5b5b",x"83d00a5c",x"78087081",x"06515271",x"9d389c84",x"085372f0",x"389c8008",x"5287e872",x"27e63872",x"7e0c7283",x"900a0c98",x"a02d8290",x"0a085379",x"802e81b4",x"387280fe",x"2e098106",x"80f43876",x"802ec138",x"807d7857",x"575a8277",x"27ffb538",x"83ffff7c",x"0c79fe18",x"53537972",x"27983880",x"dc808088",x"72555872",x"16703379",x"0c528113",x"53737326",x"f238ff15",x"76115476",x"05ff0570",x"33743370",x"72882b07",x"7f085351",x"55515271",x"732e0981",x"06feed38",x"75335372",x"8a26fee4",x"38721010",x"9af40576",x"52700851",x"52712dfe",x"d3397280",x"fd2e0981",x"06863881",x"5bfec539",x"76829f26",x"9e387a80",x"2e873880",x"73a03254",x"5b80d73d",x"7705fde0",x"05527272",x"34811757",x"fea23980",x"5afe9d39",x"7280fe2e",x"098106fe",x"93387957",x"ff7c0c81",x"775c5afe",x"8739ff3d",x"0d735280",x"5194d92d",x"833d0d04",x"81fff80d",x"8cfd0481",x"fff80da0",x"88048808",x"80c08080",x"8808a080",x"082d5088",x"0c810b90",x"0a0c0480",x"700cfaad",x"95b4da0b",x"81808071",x"710c7180",x"082e8738",x"70115198",x"cf045198",x"922dfb3d",x"0d777955",x"55805675",x"7524ab38",x"8074249d",x"38805373",x"52745180",x"e13f8808",x"5475802e",x"85388808",x"30547388",x"0c873d0d",x"04733076",x"81325754",x"dc397430",x"55815673",x"8025d238",x"ec39fa3d",x"0d787a57",x"55805776",x"7524a438",x"759f2c54",x"81537574",x"32743152",x"74519b3f",x"88085476",x"802e8538",x"88083054",x"73880c88",x"3d0d0474",x"30558157",x"d739fc3d",x"0d767853",x"54815380",x"74732652",x"5572802e",x"98387080",x"2ea93880",x"7224a438",x"71107310",x"75722653",x"545272ea",x"38735178",x"83387451",x"70880c86",x"3d0d0472",x"812a7281",x"2a535372",x"802ee638",x"717426ef",x"38737231",x"75740774",x"812a7481",x"2a555556",x"54e539ff",x"3d0d9c90",x"0bfc0570",x"08525270",x"ff2e9138",x"702dfc12",x"70085252",x"70ff2e09",x"8106f138",x"833d0d04",x"04eebc3f",x"04000000",x"00ffffff",x"ff00ffff",x"ffff00ff",x"ffffff00",x"00000964",x"00000996",x"0000093e",x"000007c9",x"000009ed",x"00000a04",x"0000085c",x"000008eb",x"00000775",x"00000a18",x"43500d0a",x"00000000",x"4c6f6164",x"65642c20",x"73746172",x"74696e67",x"2e2e2e0d",x"0a000000",x"0d0a5a50",x"55494e4f",x"0d0a0000",x"00000000",x"00000000",x"00000000",x"00000e18",x"01090460",x"00000000",x"05b8d800",x"b4010f00",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"ffffffff",x"00000000",x"ffffffff",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000");

begin

  process (clk)
  begin
    if rising_edge(clk) then
      if ENA='1' then
        if WEA='1' then
          RAM(conv_integer(ADDRA) ) := DIA;
        end if;
        DOA <= RAM(conv_integer(ADDRA)) ;
      end if;
    end if;
  end process;  

  process (clk)
  begin
    if rising_edge(clk) then
      if ENB='1' then
        if WEB='1' then
          RAM( conv_integer(ADDRB) ) := DIB;
        end if;
        DOB <= RAM(conv_integer(ADDRB)) ;
      end if;
    end if;
  end process;  
end behave;
