library IEEE;
use IEEE.std_logic_1164.all; 
use IEEE.std_logic_unsigned.all; 
use ieee.numeric_std.all;

entity bootloader_dp_32 is
  port (
    CLK:              in std_logic;
    WEA:  in std_logic;
    ENA:  in std_logic;
    MASKA:    in std_logic_vector(3 downto 0);
    ADDRA:         in std_logic_vector(11 downto 2);
    DIA:        in std_logic_vector(31 downto 0);
    DOA:         out std_logic_vector(31 downto 0);
    WEB:  in std_logic;
    ENB:  in std_logic;
    ADDRB:         in std_logic_vector(11 downto 2);
    DIB:        in std_logic_vector(31 downto 0);
    MASKB:    in std_logic_vector(3 downto 0);
    DOB:         out std_logic_vector(31 downto 0)
  );
end entity bootloader_dp_32;

architecture behave of bootloader_dp_32 is

  subtype RAM_WORD is STD_LOGIC_VECTOR (31 downto 0);
  type RAM_TABLE is array (0 to 1023) of RAM_WORD;
 shared variable RAM: RAM_TABLE := RAM_TABLE'(
x"0b0b0b97",x"f2040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b97",x"d3040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fd0608",x"72830609",x"81058205",x"832b2a83",x"ffff0652",x"04000000",x"00000000",x"00000000",x"71fd0608",x"83ffff73",x"83060981",x"05820583",x"2b2b0906",x"7383ffff",x"0b0b0b0b",x"83a70400",x"72098105",x"72057373",x"09060906",x"73097306",x"070a8106",x"53510400",x"00000000",x"00000000",x"72722473",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71737109",x"71068106",x"30720a10",x"0a720a10",x"0a31050a",x"81065151",x"53510400",x"00000000",x"72722673",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"cc040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"720a722b",x"0a535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72729f06",x"0981050b",x"0b0b88af",x"05040000",x"00000000",x"00000000",x"00000000",x"00000000",x"72722aff",x"739f062a",x"0974090a",x"8106ff05",x"06075351",x"04000000",x"00000000",x"00000000",x"71715351",x"020d0406",x"73830609",x"81058205",x"832b0b2b",x"0772fc06",x"0c515104",x"00000000",x"72098105",x"72050970",x"81050906",x"0a810653",x"51040000",x"00000000",x"00000000",x"00000000",x"72098105",x"72050970",x"81050906",x"0a098106",x"53510400",x"00000000",x"00000000",x"00000000",x"71098105",x"52040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72720981",x"05055351",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097206",x"73730906",x"07535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fc0608",x"72830609",x"81058305",x"1010102a",x"81ff0652",x"04000000",x"00000000",x"00000000",x"71fc0608",x"0b0b0b9e",x"9c738306",x"10100508",x"060b0b0b",x"88b20400",x"00000000",x"00000000",x"0b0b0b89",x"80040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"e8040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097081",x"0509060a",x"8106ff05",x"70547106",x"73097274",x"05ff0506",x"07515151",x"04000000",x"72097081",x"0509060a",x"098106ff",x"05705471",x"06730972",x"7405ff05",x"06075151",x"51040000",x"05ff0504",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"810b0b0b",x"0b9f940c",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71810552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"02840572",x"10100552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"717105ff",x"05715351",x"020d0400",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"81dd3f95",x"ea3f0400",x"00000000",x"00000000",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101053",x"51047381",x"ff067383",x"06098105",x"83051010",x"102b0772",x"fc060c51",x"51043c04",x"72728072",x"8106ff05",x"09720605",x"71105272",x"0a100a53",x"72ed3851",x"51535104",x"88088c08",x"90087575",x"999d2d50",x"50880856",x"900c8c0c",x"880c5104",x"88088c08",x"90087575",x"98d92d50",x"50880856",x"900c8c0c",x"880c5104",x"88088c08",x"90088ebb",x"2d900c8c",x"0c880c04",x"ff3d0d0b",x"0b0b9fa4",x"335170a6",x"389fa008",x"70085252",x"70802e92",x"3884129f",x"a00c702d",x"9fa00870",x"08525270",x"f038810b",x"0b0b0b9f",x"a434833d",x"0d040480",x"3d0d0b0b",x"0b9fd008",x"802e8e38",x"0b0b0b0b",x"800b802e",x"09810685",x"38823d0d",x"040b0b0b",x"9fd0510b",x"0b0bf5f8",x"3f823d0d",x"0404ff3d",x"0d80c480",x"80845271",x"0870822a",x"70810651",x"515170f3",x"38833d0d",x"04ff3d0d",x"80c48080",x"84527108",x"70812a70",x"81065151",x"5170f338",x"7382900a",x"0c833d0d",x"04fd3d0d",x"75547333",x"7081ff06",x"53537180",x"2e8e3872",x"81ff0651",x"8aa92d81",x"1454e739",x"853d0d04",x"fe3d0d74",x"7080dc80",x"80880c70",x"81ff06ff",x"83115451",x"53718126",x"8d3880fd",x"518aa92d",x"72a03251",x"83397251",x"8aa92d84",x"3d0d0480",x"3d0d83ff",x"ff0b83d0",x"0a0c80fe",x"518aa92d",x"823d0d04",x"ff3d0d83",x"d00a0870",x"882a5252",x"8aec2d71",x"81ff0651",x"8aec2d80",x"fe518aa9",x"2d833d0d",x"0482f6ff",x"0b80cc80",x"80880c80",x"0b80cc80",x"80840c9f",x"0b83900a",x"0c04ff3d",x"0d737008",x"515180c8",x"80808470",x"08708480",x"8007720c",x"5252833d",x"0d04ff3d",x"0d80c880",x"80847008",x"70fbffff",x"06720c52",x"52833d0d",x"04a0900b",x"a0800c9f",x"a80ba084",x"0c988b2d",x"ff3d0d73",x"518b710c",x"90115298",x"8080720c",x"80720c70",x"0883ffff",x"06880c83",x"3d0d04fa",x"3d0d787a",x"7dff1e57",x"57585373",x"ff2ea738",x"80568452",x"75730c72",x"0888180c",x"ff125271",x"f3387484",x"16740872",x"0cff1656",x"565273ff",x"2e098106",x"dd38883d",x"0d04f83d",x"0d80c080",x"80845783",x"d00a0b9e",x"e452598a",x"c92d8c86",x"2d76518c",x"ac2d9fa8",x"70880810",x"10988084",x"05717084",x"05530c56",x"56fb8084",x"a1ad750c",x"9ed40b88",x"170c8070",x"780c770c",x"760883ff",x"ff065683",x"ffdf800b",x"8808278f",x"389eec51",x"8ac92d9f",x"90518ac9",x"2dff3983",x"ffff790c",x"a0805488",x"08537852",x"76518ccb",x"2d76518b",x"ea2d7808",x"5574762e",x"893880c3",x"518aa92d",x"ff39a084",x"085574fa",x"a090ae80",x"2e893880",x"c2518aa9",x"2dff399e",x"f0518ac9",x"2d900a70",x"0870ffbf",x"06720c56",x"568a8e2d",x"8c9d2dff",x"3d0d9fb4",x"0881119f",x"b40c5183",x"900a7008",x"70feff06",x"720c5252",x"833d0d04",x"803d0d8b",x"9b2d7281",x"8007518a",x"ec2d8bb0",x"2d823d0d",x"04fe3d0d",x"80c08080",x"84538c86",x"2d85730c",x"80730c72",x"087081ff",x"06745351",x"528bea2d",x"71880c84",x"3d0d0404",x"f93d0d79",x"5780c080",x"8084568c",x"862d8117",x"33821833",x"71828029",x"05535371",x"802e9438",x"85177255",x"53727081",x"05543376",x"0cff1454",x"73f33883",x"17338418",x"33718280",x"29055652",x"80547375",x"27973873",x"5877760c",x"73177608",x"53537173",x"34811454",x"747426ed",x"3875518b",x"ea2d8b9b",x"2d818451",x"8aec2d74",x"882a518a",x"ec2d7451",x"8aec2d80",x"54737527",x"8f387317",x"70335252",x"8aec2d81",x"1454ee39",x"8bb02d89",x"3d0d04f9",x"3d0d7956",x"80c08080",x"84558c86",x"2d86750c",x"74518bea",x"2d8c862d",x"81ad7076",x"0c811733",x"82183371",x"82802905",x"83193378",x"0c841933",x"780c8519",x"33780c59",x"53538054",x"737727b3",x"38725873",x"802e8738",x"8c862d77",x"750c7316",x"86113376",x"0c871133",x"760c5274",x"518bea2d",x"8eed2d88",x"08810652",x"71f63882",x"14547674",x"26d1388c",x"862d8475",x"0c74518b",x"ea2d8b9b",x"2d818751",x"8aec2d8b",x"b02d893d",x"0d04fc3d",x"0d768111",x"33821233",x"71902b71",x"882b0783",x"14337072",x"07882b84",x"16337107",x"51525357",x"57545288",x"518ed82d",x"81ff518a",x"a92d80c4",x"80808453",x"72087081",x"2a708106",x"51515271",x"f3387384",x"80800780",x"c4808084",x"0c863d0d",x"04fe3d0d",x"8eed2d88",x"08880881",x"06535371",x"f3388b9b",x"2d818351",x"8aec2d72",x"518aec2d",x"8bb02d84",x"3d0d04fe",x"3d0d800b",x"9fb40c8b",x"9b2d8181",x"518aec2d",x"9ed4538f",x"52727081",x"05543351",x"8aec2dff",x"125271ff",x"2e098106",x"ec388bb0",x"2d843d0d",x"04fe3d0d",x"800b9fb4",x"0c8b9b2d",x"8182518a",x"ec2d80c0",x"80808452",x"8c862d81",x"f90a0b80",x"c080809c",x"0c710872",x"52538bea",x"2d729fbc",x"0c72902a",x"518aec2d",x"9fbc0888",x"2a518aec",x"2d9fbc08",x"518aec2d",x"8eed2d88",x"08518aec",x"2d8bb02d",x"843d0d04",x"803d0d81",x"0b9fb80c",x"800b8390",x"0a0c8551",x"8ed82d82",x"3d0d0480",x"3d0d800b",x"9fb80c8b",x"d12d8651",x"8ed82d82",x"3d0d04fd",x"3d0d80c0",x"80808454",x"8a518ed8",x"2d8c862d",x"9fa87452",x"538cac2d",x"72880810",x"10988084",x"05717084",x"05530c52",x"fb8084a1",x"ad720c9e",x"d40b8814",x"0c73518b",x"ea2d8a8e",x"2d8c9d2d",x"ffab3d0d",x"800b9fb8",x"0c800b9f",x"b40c800b",x"8ebb0ba0",x"800c5780",x"c4808084",x"558480b3",x"750c80c8",x"8080a453",x"fbffff73",x"08707206",x"750c5354",x"80c88080",x"94700870",x"7606720c",x"5353a870",x"99d57170",x"8405530c",x"9ab2710c",x"539bcb0b",x"88120c9c",x"da0b8c12",x"0c53880b",x"80d08080",x"840c80d0",x"0a538173",x"0c9f8851",x"8ac92d8b",x"d12d8288",x"880b80dc",x"8080840c",x"81f20b90",x"0a0c80c0",x"80808470",x"52528bea",x"2d8c862d",x"71518bea",x"2d8c862d",x"84720c71",x"518bea2d",x"76777675",x"933d4141",x"5b5b5b83",x"d00a5c78",x"08708106",x"5152719d",x"389fb808",x"5372f038",x"9fb40852",x"87e87227",x"e638727e",x"0c728390",x"0a0c9883",x"2d82900a",x"08537980",x"2e81b438",x"7280fe2e",x"09810680",x"f4387680",x"2ec13880",x"7d785856",x"5a827727",x"ffb53883",x"ffff7c0c",x"79fe1853",x"53797227",x"983880dc",x"80808872",x"55587215",x"7033790c",x"52811353",x"737326f2",x"38ff1675",x"11547505",x"ff057033",x"74337072",x"882b077f",x"08535155",x"51527173",x"2e098106",x"feed3874",x"3353728a",x"26fee438",x"7210109e",x"a8057552",x"70085152",x"712dfed3",x"397280fd",x"2e098106",x"8638815b",x"fec53976",x"829f269e",x"387a802e",x"87388073",x"a032545b",x"80d73d77",x"05fde005",x"52727234",x"811757fe",x"a239805a",x"fe9d3972",x"80fe2e09",x"8106fe93",x"38795783",x"ffff7c0c",x"81775c5a",x"fe853980",x"3d0d8808",x"8c089008",x"a0800851",x"702d900c",x"8c0c8a0c",x"810b80d0",x"0a0c823d",x"0d04ff3d",x"0d98ad2d",x"80528051",x"94a42d83",x"3d0d0483",x"fffff80d",x"8d860483",x"fffff80d",x"a0880400",x"00000000",x"00000000",x"00000000",x"820b80d0",x"8080900c",x"0b0b0b04",x"0083f00a",x"0b800ba0",x"80721208",x"720c8412",x"5271712e",x"ff05f238",x"028c050d",x"98a00400",x"00000000",x"00000000",x"00000000",x"00fb3d0d",x"77795555",x"80567575",x"24ab3880",x"74249d38",x"80537352",x"745180e1",x"3f880854",x"75802e85",x"38880830",x"5473880c",x"873d0d04",x"73307681",x"325754dc",x"39743055",x"81567380",x"25d238ec",x"39fa3d0d",x"787a5755",x"80577675",x"24a43875",x"9f2c5481",x"53757432",x"74315274",x"519b3f88",x"08547680",x"2e853888",x"08305473",x"880c883d",x"0d047430",x"558157d7",x"39fc3d0d",x"76785354",x"81538074",x"73265255",x"72802e98",x"3870802e",x"a9388072",x"24a43871",x"10731075",x"72265354",x"5272ea38",x"73517883",x"38745170",x"880c863d",x"0d047281",x"2a72812a",x"53537280",x"2ee63871",x"7426ef38",x"73723175",x"74077481",x"2a74812a",x"55555654",x"e539fc3d",x"0d767079",x"7b555555",x"558f7227",x"8c387275",x"07830651",x"70802ea7",x"38ff1252",x"71ff2e98",x"38727081",x"05543374",x"70810556",x"34ff1252",x"71ff2e09",x"8106ea38",x"74880c86",x"3d0d0474",x"51727084",x"05540871",x"70840553",x"0c727084",x"05540871",x"70840553",x"0c727084",x"05540871",x"70840553",x"0c727084",x"05540871",x"70840553",x"0cf01252",x"718f26c9",x"38837227",x"95387270",x"84055408",x"71708405",x"530cfc12",x"52718326",x"ed387054",x"ff8339fc",x"3d0d7679",x"71028c05",x"9f053357",x"55535583",x"72278a38",x"74830651",x"70802ea2",x"38ff1252",x"71ff2e93",x"38737370",x"81055534",x"ff125271",x"ff2e0981",x"06ef3874",x"880c863d",x"0d047474",x"882b7507",x"7071902b",x"07515451",x"8f7227a5",x"38727170",x"8405530c",x"72717084",x"05530c72",x"71708405",x"530c7271",x"70840553",x"0cf01252",x"718f26dd",x"38837227",x"90387271",x"70840553",x"0cfc1252",x"718326f2",x"387053ff",x"9039fb3d",x"0d777970",x"72078306",x"53545270",x"93387173",x"73085456",x"54717308",x"2e80c438",x"73755452",x"71337081",x"ff065254",x"70802e9d",x"38723355",x"70752e09",x"81069538",x"81128114",x"71337081",x"ff065456",x"545270e5",x"38723355",x"7381ff06",x"7581ff06",x"71713188",x"0c525287",x"3d0d0471",x"0970f7fb",x"fdff1406",x"70f88482",x"81800651",x"51517097",x"38841484",x"16710854",x"56547175",x"082edc38",x"73755452",x"ff963980",x"0b880c87",x"3d0d04ff",x"3d0d9fc4",x"0bfc0570",x"08525270",x"ff2e9138",x"702dfc12",x"70085252",x"70ff2e09",x"8106f138",x"833d0d04",x"04eb913f",x"04000000",x"00ffffff",x"ff00ffff",x"ffff00ff",x"ffffff00",x"0000092f",x"00000961",x"00000909",x"00000794",x"000009b8",x"000009cf",x"00000827",x"000008b6",x"00000793",x"000009e3",x"01090600",x"007fef80",x"05b8d800",x"a4041700",x"43500d0a",x"00000000",x"534c4b00",x"4c6f6164",x"65642c20",x"73746172",x"74696e67",x"2e2e2e0d",x"0a000000",x"0d0a5a50",x"55494e4f",x"0d0a0000",x"00000000",x"00000000",x"00000000",x"00000fcc",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"ffffffff",x"00000000",x"ffffffff",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000");

begin

  process (clk)
  begin
    if rising_edge(clk) then
      if ENA='1' then
        if WEA='1' then
          RAM(conv_integer(ADDRA) ) := DIA;
        end if;
        DOA <= RAM(conv_integer(ADDRA)) ;
      end if;
    end if;
  end process;  

  process (clk)
  begin
    if rising_edge(clk) then
      if ENB='1' then
        if WEB='1' then
          RAM( conv_integer(ADDRB) ) := DIB;
        end if;
        DOB <= RAM(conv_integer(ADDRB)) ;
      end if;
    end if;
  end process;  
end behave;
