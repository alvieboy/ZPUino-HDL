---------------------------------------------------------------------
--	Filename:	gh_sincos_rom_16_2.vhd
--			
--	Description:
--		Sin Cos look up table 16 bit (from 1/2 table)
--
--	Copyright (c) 2008 by George Huber 
--		an OpenCores.org Project
--		free to use, but see documentation for conditions 
--
--	Revision 	History:
--	Revision 	Date      	Author   	Comment
--	-------- 	----------	---------	-----------
--	1.0      	10/26/08  	h LeFevre	Initial revision
--	
------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

entity gh_sincos_rom_16_2 is
	port (
		CLK : in std_logic;
		ADD : in std_logic_vector(15 downto 0);
		sin : out std_logic_vector(15 downto 0);
		cos : out std_logic_vector(15 downto 0)
		);
end entity;

architecture a of gh_sincos_rom_16_2 is

	signal dADD :  STD_LOGIC;
	signal msin, mcos :  STD_LOGIC_VECTOR(15 DOWNTO 0);

	type rom_mem is array (0 to 32767) of std_logic_vector (15 downto 0);
	constant isin : rom_mem :=(  
    x"0000", x"0003", x"0006", x"0009", x"000d", x"0010", x"0013", x"0016", 
    x"0019", x"001c", x"001f", x"0023", x"0026", x"0029", x"002c", x"002f", 
    x"0032", x"0035", x"0039", x"003c", x"003f", x"0042", x"0045", x"0048", 
    x"004b", x"004f", x"0052", x"0055", x"0058", x"005b", x"005e", x"0061", 
    x"0065", x"0068", x"006b", x"006e", x"0071", x"0074", x"0077", x"007b", 
    x"007e", x"0081", x"0084", x"0087", x"008a", x"008d", x"0091", x"0094", 
    x"0097", x"009a", x"009d", x"00a0", x"00a3", x"00a6", x"00aa", x"00ad", 
    x"00b0", x"00b3", x"00b6", x"00b9", x"00bc", x"00c0", x"00c3", x"00c6", 
    x"00c9", x"00cc", x"00cf", x"00d2", x"00d6", x"00d9", x"00dc", x"00df", 
    x"00e2", x"00e5", x"00e8", x"00ec", x"00ef", x"00f2", x"00f5", x"00f8", 
    x"00fb", x"00fe", x"0102", x"0105", x"0108", x"010b", x"010e", x"0111", 
    x"0114", x"0118", x"011b", x"011e", x"0121", x"0124", x"0127", x"012a", 
    x"012e", x"0131", x"0134", x"0137", x"013a", x"013d", x"0140", x"0144", 
    x"0147", x"014a", x"014d", x"0150", x"0153", x"0156", x"015a", x"015d", 
    x"0160", x"0163", x"0166", x"0169", x"016c", x"0170", x"0173", x"0176", 
    x"0179", x"017c", x"017f", x"0182", x"0186", x"0189", x"018c", x"018f", 
    x"0192", x"0195", x"0198", x"019c", x"019f", x"01a2", x"01a5", x"01a8", 
    x"01ab", x"01ae", x"01b2", x"01b5", x"01b8", x"01bb", x"01be", x"01c1", 
    x"01c4", x"01c8", x"01cb", x"01ce", x"01d1", x"01d4", x"01d7", x"01da", 
    x"01dd", x"01e1", x"01e4", x"01e7", x"01ea", x"01ed", x"01f0", x"01f3", 
    x"01f7", x"01fa", x"01fd", x"0200", x"0203", x"0206", x"0209", x"020d", 
    x"0210", x"0213", x"0216", x"0219", x"021c", x"021f", x"0223", x"0226", 
    x"0229", x"022c", x"022f", x"0232", x"0235", x"0239", x"023c", x"023f", 
    x"0242", x"0245", x"0248", x"024b", x"024f", x"0252", x"0255", x"0258", 
    x"025b", x"025e", x"0261", x"0265", x"0268", x"026b", x"026e", x"0271", 
    x"0274", x"0277", x"027b", x"027e", x"0281", x"0284", x"0287", x"028a", 
    x"028d", x"0291", x"0294", x"0297", x"029a", x"029d", x"02a0", x"02a3", 
    x"02a7", x"02aa", x"02ad", x"02b0", x"02b3", x"02b6", x"02b9", x"02bd", 
    x"02c0", x"02c3", x"02c6", x"02c9", x"02cc", x"02cf", x"02d2", x"02d6", 
    x"02d9", x"02dc", x"02df", x"02e2", x"02e5", x"02e8", x"02ec", x"02ef", 
    x"02f2", x"02f5", x"02f8", x"02fb", x"02fe", x"0302", x"0305", x"0308", 
    x"030b", x"030e", x"0311", x"0314", x"0318", x"031b", x"031e", x"0321", 
    x"0324", x"0327", x"032a", x"032e", x"0331", x"0334", x"0337", x"033a", 
    x"033d", x"0340", x"0344", x"0347", x"034a", x"034d", x"0350", x"0353", 
    x"0356", x"035a", x"035d", x"0360", x"0363", x"0366", x"0369", x"036c", 
    x"0370", x"0373", x"0376", x"0379", x"037c", x"037f", x"0382", x"0385", 
    x"0389", x"038c", x"038f", x"0392", x"0395", x"0398", x"039b", x"039f", 
    x"03a2", x"03a5", x"03a8", x"03ab", x"03ae", x"03b1", x"03b5", x"03b8", 
    x"03bb", x"03be", x"03c1", x"03c4", x"03c7", x"03cb", x"03ce", x"03d1", 
    x"03d4", x"03d7", x"03da", x"03dd", x"03e1", x"03e4", x"03e7", x"03ea", 
    x"03ed", x"03f0", x"03f3", x"03f7", x"03fa", x"03fd", x"0400", x"0403", 
    x"0406", x"0409", x"040d", x"0410", x"0413", x"0416", x"0419", x"041c", 
    x"041f", x"0423", x"0426", x"0429", x"042c", x"042f", x"0432", x"0435", 
    x"0438", x"043c", x"043f", x"0442", x"0445", x"0448", x"044b", x"044e", 
    x"0452", x"0455", x"0458", x"045b", x"045e", x"0461", x"0464", x"0468", 
    x"046b", x"046e", x"0471", x"0474", x"0477", x"047a", x"047e", x"0481", 
    x"0484", x"0487", x"048a", x"048d", x"0490", x"0494", x"0497", x"049a", 
    x"049d", x"04a0", x"04a3", x"04a6", x"04aa", x"04ad", x"04b0", x"04b3", 
    x"04b6", x"04b9", x"04bc", x"04bf", x"04c3", x"04c6", x"04c9", x"04cc", 
    x"04cf", x"04d2", x"04d5", x"04d9", x"04dc", x"04df", x"04e2", x"04e5", 
    x"04e8", x"04eb", x"04ef", x"04f2", x"04f5", x"04f8", x"04fb", x"04fe", 
    x"0501", x"0505", x"0508", x"050b", x"050e", x"0511", x"0514", x"0517", 
    x"051b", x"051e", x"0521", x"0524", x"0527", x"052a", x"052d", x"0530", 
    x"0534", x"0537", x"053a", x"053d", x"0540", x"0543", x"0546", x"054a", 
    x"054d", x"0550", x"0553", x"0556", x"0559", x"055c", x"0560", x"0563", 
    x"0566", x"0569", x"056c", x"056f", x"0572", x"0576", x"0579", x"057c", 
    x"057f", x"0582", x"0585", x"0588", x"058c", x"058f", x"0592", x"0595", 
    x"0598", x"059b", x"059e", x"05a1", x"05a5", x"05a8", x"05ab", x"05ae", 
    x"05b1", x"05b4", x"05b7", x"05bb", x"05be", x"05c1", x"05c4", x"05c7", 
    x"05ca", x"05cd", x"05d1", x"05d4", x"05d7", x"05da", x"05dd", x"05e0", 
    x"05e3", x"05e7", x"05ea", x"05ed", x"05f0", x"05f3", x"05f6", x"05f9", 
    x"05fc", x"0600", x"0603", x"0606", x"0609", x"060c", x"060f", x"0612", 
    x"0616", x"0619", x"061c", x"061f", x"0622", x"0625", x"0628", x"062c", 
    x"062f", x"0632", x"0635", x"0638", x"063b", x"063e", x"0642", x"0645", 
    x"0648", x"064b", x"064e", x"0651", x"0654", x"0657", x"065b", x"065e", 
    x"0661", x"0664", x"0667", x"066a", x"066d", x"0671", x"0674", x"0677", 
    x"067a", x"067d", x"0680", x"0683", x"0687", x"068a", x"068d", x"0690", 
    x"0693", x"0696", x"0699", x"069d", x"06a0", x"06a3", x"06a6", x"06a9", 
    x"06ac", x"06af", x"06b2", x"06b6", x"06b9", x"06bc", x"06bf", x"06c2", 
    x"06c5", x"06c8", x"06cc", x"06cf", x"06d2", x"06d5", x"06d8", x"06db", 
    x"06de", x"06e2", x"06e5", x"06e8", x"06eb", x"06ee", x"06f1", x"06f4", 
    x"06f7", x"06fb", x"06fe", x"0701", x"0704", x"0707", x"070a", x"070d", 
    x"0711", x"0714", x"0717", x"071a", x"071d", x"0720", x"0723", x"0727", 
    x"072a", x"072d", x"0730", x"0733", x"0736", x"0739", x"073c", x"0740", 
    x"0743", x"0746", x"0749", x"074c", x"074f", x"0752", x"0756", x"0759", 
    x"075c", x"075f", x"0762", x"0765", x"0768", x"076c", x"076f", x"0772", 
    x"0775", x"0778", x"077b", x"077e", x"0781", x"0785", x"0788", x"078b", 
    x"078e", x"0791", x"0794", x"0797", x"079b", x"079e", x"07a1", x"07a4", 
    x"07a7", x"07aa", x"07ad", x"07b1", x"07b4", x"07b7", x"07ba", x"07bd", 
    x"07c0", x"07c3", x"07c6", x"07ca", x"07cd", x"07d0", x"07d3", x"07d6", 
    x"07d9", x"07dc", x"07e0", x"07e3", x"07e6", x"07e9", x"07ec", x"07ef", 
    x"07f2", x"07f6", x"07f9", x"07fc", x"07ff", x"0802", x"0805", x"0808", 
    x"080b", x"080f", x"0812", x"0815", x"0818", x"081b", x"081e", x"0821", 
    x"0825", x"0828", x"082b", x"082e", x"0831", x"0834", x"0837", x"083a", 
    x"083e", x"0841", x"0844", x"0847", x"084a", x"084d", x"0850", x"0854", 
    x"0857", x"085a", x"085d", x"0860", x"0863", x"0866", x"086a", x"086d", 
    x"0870", x"0873", x"0876", x"0879", x"087c", x"087f", x"0883", x"0886", 
    x"0889", x"088c", x"088f", x"0892", x"0895", x"0899", x"089c", x"089f", 
    x"08a2", x"08a5", x"08a8", x"08ab", x"08ae", x"08b2", x"08b5", x"08b8", 
    x"08bb", x"08be", x"08c1", x"08c4", x"08c8", x"08cb", x"08ce", x"08d1", 
    x"08d4", x"08d7", x"08da", x"08dd", x"08e1", x"08e4", x"08e7", x"08ea", 
    x"08ed", x"08f0", x"08f3", x"08f7", x"08fa", x"08fd", x"0900", x"0903", 
    x"0906", x"0909", x"090c", x"0910", x"0913", x"0916", x"0919", x"091c", 
    x"091f", x"0922", x"0926", x"0929", x"092c", x"092f", x"0932", x"0935", 
    x"0938", x"093b", x"093f", x"0942", x"0945", x"0948", x"094b", x"094e", 
    x"0951", x"0955", x"0958", x"095b", x"095e", x"0961", x"0964", x"0967", 
    x"096a", x"096e", x"0971", x"0974", x"0977", x"097a", x"097d", x"0980", 
    x"0984", x"0987", x"098a", x"098d", x"0990", x"0993", x"0996", x"0999", 
    x"099d", x"09a0", x"09a3", x"09a6", x"09a9", x"09ac", x"09af", x"09b3", 
    x"09b6", x"09b9", x"09bc", x"09bf", x"09c2", x"09c5", x"09c8", x"09cc", 
    x"09cf", x"09d2", x"09d5", x"09d8", x"09db", x"09de", x"09e2", x"09e5", 
    x"09e8", x"09eb", x"09ee", x"09f1", x"09f4", x"09f7", x"09fb", x"09fe", 
    x"0a01", x"0a04", x"0a07", x"0a0a", x"0a0d", x"0a11", x"0a14", x"0a17", 
    x"0a1a", x"0a1d", x"0a20", x"0a23", x"0a26", x"0a2a", x"0a2d", x"0a30", 
    x"0a33", x"0a36", x"0a39", x"0a3c", x"0a3f", x"0a43", x"0a46", x"0a49", 
    x"0a4c", x"0a4f", x"0a52", x"0a55", x"0a59", x"0a5c", x"0a5f", x"0a62", 
    x"0a65", x"0a68", x"0a6b", x"0a6e", x"0a72", x"0a75", x"0a78", x"0a7b", 
    x"0a7e", x"0a81", x"0a84", x"0a87", x"0a8b", x"0a8e", x"0a91", x"0a94", 
    x"0a97", x"0a9a", x"0a9d", x"0aa1", x"0aa4", x"0aa7", x"0aaa", x"0aad", 
    x"0ab0", x"0ab3", x"0ab6", x"0aba", x"0abd", x"0ac0", x"0ac3", x"0ac6", 
    x"0ac9", x"0acc", x"0acf", x"0ad3", x"0ad6", x"0ad9", x"0adc", x"0adf", 
    x"0ae2", x"0ae5", x"0ae9", x"0aec", x"0aef", x"0af2", x"0af5", x"0af8", 
    x"0afb", x"0afe", x"0b02", x"0b05", x"0b08", x"0b0b", x"0b0e", x"0b11", 
    x"0b14", x"0b17", x"0b1b", x"0b1e", x"0b21", x"0b24", x"0b27", x"0b2a", 
    x"0b2d", x"0b31", x"0b34", x"0b37", x"0b3a", x"0b3d", x"0b40", x"0b43", 
    x"0b46", x"0b4a", x"0b4d", x"0b50", x"0b53", x"0b56", x"0b59", x"0b5c", 
    x"0b5f", x"0b63", x"0b66", x"0b69", x"0b6c", x"0b6f", x"0b72", x"0b75", 
    x"0b78", x"0b7c", x"0b7f", x"0b82", x"0b85", x"0b88", x"0b8b", x"0b8e", 
    x"0b92", x"0b95", x"0b98", x"0b9b", x"0b9e", x"0ba1", x"0ba4", x"0ba7", 
    x"0bab", x"0bae", x"0bb1", x"0bb4", x"0bb7", x"0bba", x"0bbd", x"0bc0", 
    x"0bc4", x"0bc7", x"0bca", x"0bcd", x"0bd0", x"0bd3", x"0bd6", x"0bd9", 
    x"0bdd", x"0be0", x"0be3", x"0be6", x"0be9", x"0bec", x"0bef", x"0bf3", 
    x"0bf6", x"0bf9", x"0bfc", x"0bff", x"0c02", x"0c05", x"0c08", x"0c0c", 
    x"0c0f", x"0c12", x"0c15", x"0c18", x"0c1b", x"0c1e", x"0c21", x"0c25", 
    x"0c28", x"0c2b", x"0c2e", x"0c31", x"0c34", x"0c37", x"0c3a", x"0c3e", 
    x"0c41", x"0c44", x"0c47", x"0c4a", x"0c4d", x"0c50", x"0c53", x"0c57", 
    x"0c5a", x"0c5d", x"0c60", x"0c63", x"0c66", x"0c69", x"0c6c", x"0c70", 
    x"0c73", x"0c76", x"0c79", x"0c7c", x"0c7f", x"0c82", x"0c85", x"0c89", 
    x"0c8c", x"0c8f", x"0c92", x"0c95", x"0c98", x"0c9b", x"0c9e", x"0ca2", 
    x"0ca5", x"0ca8", x"0cab", x"0cae", x"0cb1", x"0cb4", x"0cb7", x"0cbb", 
    x"0cbe", x"0cc1", x"0cc4", x"0cc7", x"0cca", x"0ccd", x"0cd1", x"0cd4", 
    x"0cd7", x"0cda", x"0cdd", x"0ce0", x"0ce3", x"0ce6", x"0cea", x"0ced", 
    x"0cf0", x"0cf3", x"0cf6", x"0cf9", x"0cfc", x"0cff", x"0d03", x"0d06", 
    x"0d09", x"0d0c", x"0d0f", x"0d12", x"0d15", x"0d18", x"0d1c", x"0d1f", 
    x"0d22", x"0d25", x"0d28", x"0d2b", x"0d2e", x"0d31", x"0d35", x"0d38", 
    x"0d3b", x"0d3e", x"0d41", x"0d44", x"0d47", x"0d4a", x"0d4e", x"0d51", 
    x"0d54", x"0d57", x"0d5a", x"0d5d", x"0d60", x"0d63", x"0d66", x"0d6a", 
    x"0d6d", x"0d70", x"0d73", x"0d76", x"0d79", x"0d7c", x"0d7f", x"0d83", 
    x"0d86", x"0d89", x"0d8c", x"0d8f", x"0d92", x"0d95", x"0d98", x"0d9c", 
    x"0d9f", x"0da2", x"0da5", x"0da8", x"0dab", x"0dae", x"0db1", x"0db5", 
    x"0db8", x"0dbb", x"0dbe", x"0dc1", x"0dc4", x"0dc7", x"0dca", x"0dce", 
    x"0dd1", x"0dd4", x"0dd7", x"0dda", x"0ddd", x"0de0", x"0de3", x"0de7", 
    x"0dea", x"0ded", x"0df0", x"0df3", x"0df6", x"0df9", x"0dfc", x"0e00", 
    x"0e03", x"0e06", x"0e09", x"0e0c", x"0e0f", x"0e12", x"0e15", x"0e19", 
    x"0e1c", x"0e1f", x"0e22", x"0e25", x"0e28", x"0e2b", x"0e2e", x"0e32", 
    x"0e35", x"0e38", x"0e3b", x"0e3e", x"0e41", x"0e44", x"0e47", x"0e4a", 
    x"0e4e", x"0e51", x"0e54", x"0e57", x"0e5a", x"0e5d", x"0e60", x"0e63", 
    x"0e67", x"0e6a", x"0e6d", x"0e70", x"0e73", x"0e76", x"0e79", x"0e7c", 
    x"0e80", x"0e83", x"0e86", x"0e89", x"0e8c", x"0e8f", x"0e92", x"0e95", 
    x"0e99", x"0e9c", x"0e9f", x"0ea2", x"0ea5", x"0ea8", x"0eab", x"0eae", 
    x"0eb1", x"0eb5", x"0eb8", x"0ebb", x"0ebe", x"0ec1", x"0ec4", x"0ec7", 
    x"0eca", x"0ece", x"0ed1", x"0ed4", x"0ed7", x"0eda", x"0edd", x"0ee0", 
    x"0ee3", x"0ee7", x"0eea", x"0eed", x"0ef0", x"0ef3", x"0ef6", x"0ef9", 
    x"0efc", x"0eff", x"0f03", x"0f06", x"0f09", x"0f0c", x"0f0f", x"0f12", 
    x"0f15", x"0f18", x"0f1c", x"0f1f", x"0f22", x"0f25", x"0f28", x"0f2b", 
    x"0f2e", x"0f31", x"0f35", x"0f38", x"0f3b", x"0f3e", x"0f41", x"0f44", 
    x"0f47", x"0f4a", x"0f4d", x"0f51", x"0f54", x"0f57", x"0f5a", x"0f5d", 
    x"0f60", x"0f63", x"0f66", x"0f6a", x"0f6d", x"0f70", x"0f73", x"0f76", 
    x"0f79", x"0f7c", x"0f7f", x"0f82", x"0f86", x"0f89", x"0f8c", x"0f8f", 
    x"0f92", x"0f95", x"0f98", x"0f9b", x"0f9f", x"0fa2", x"0fa5", x"0fa8", 
    x"0fab", x"0fae", x"0fb1", x"0fb4", x"0fb8", x"0fbb", x"0fbe", x"0fc1", 
    x"0fc4", x"0fc7", x"0fca", x"0fcd", x"0fd0", x"0fd4", x"0fd7", x"0fda", 
    x"0fdd", x"0fe0", x"0fe3", x"0fe6", x"0fe9", x"0fec", x"0ff0", x"0ff3", 
    x"0ff6", x"0ff9", x"0ffc", x"0fff", x"1002", x"1005", x"1009", x"100c", 
    x"100f", x"1012", x"1015", x"1018", x"101b", x"101e", x"1021", x"1025", 
    x"1028", x"102b", x"102e", x"1031", x"1034", x"1037", x"103a", x"103e", 
    x"1041", x"1044", x"1047", x"104a", x"104d", x"1050", x"1053", x"1056", 
    x"105a", x"105d", x"1060", x"1063", x"1066", x"1069", x"106c", x"106f", 
    x"1072", x"1076", x"1079", x"107c", x"107f", x"1082", x"1085", x"1088", 
    x"108b", x"108f", x"1092", x"1095", x"1098", x"109b", x"109e", x"10a1", 
    x"10a4", x"10a7", x"10ab", x"10ae", x"10b1", x"10b4", x"10b7", x"10ba", 
    x"10bd", x"10c0", x"10c3", x"10c7", x"10ca", x"10cd", x"10d0", x"10d3", 
    x"10d6", x"10d9", x"10dc", x"10e0", x"10e3", x"10e6", x"10e9", x"10ec", 
    x"10ef", x"10f2", x"10f5", x"10f8", x"10fc", x"10ff", x"1102", x"1105", 
    x"1108", x"110b", x"110e", x"1111", x"1114", x"1118", x"111b", x"111e", 
    x"1121", x"1124", x"1127", x"112a", x"112d", x"1130", x"1134", x"1137", 
    x"113a", x"113d", x"1140", x"1143", x"1146", x"1149", x"114c", x"1150", 
    x"1153", x"1156", x"1159", x"115c", x"115f", x"1162", x"1165", x"1168", 
    x"116c", x"116f", x"1172", x"1175", x"1178", x"117b", x"117e", x"1181", 
    x"1185", x"1188", x"118b", x"118e", x"1191", x"1194", x"1197", x"119a", 
    x"119d", x"11a1", x"11a4", x"11a7", x"11aa", x"11ad", x"11b0", x"11b3", 
    x"11b6", x"11b9", x"11bd", x"11c0", x"11c3", x"11c6", x"11c9", x"11cc", 
    x"11cf", x"11d2", x"11d5", x"11d9", x"11dc", x"11df", x"11e2", x"11e5", 
    x"11e8", x"11eb", x"11ee", x"11f1", x"11f5", x"11f8", x"11fb", x"11fe", 
    x"1201", x"1204", x"1207", x"120a", x"120d", x"1210", x"1214", x"1217", 
    x"121a", x"121d", x"1220", x"1223", x"1226", x"1229", x"122c", x"1230", 
    x"1233", x"1236", x"1239", x"123c", x"123f", x"1242", x"1245", x"1248", 
    x"124c", x"124f", x"1252", x"1255", x"1258", x"125b", x"125e", x"1261", 
    x"1264", x"1268", x"126b", x"126e", x"1271", x"1274", x"1277", x"127a", 
    x"127d", x"1280", x"1284", x"1287", x"128a", x"128d", x"1290", x"1293", 
    x"1296", x"1299", x"129c", x"12a0", x"12a3", x"12a6", x"12a9", x"12ac", 
    x"12af", x"12b2", x"12b5", x"12b8", x"12bb", x"12bf", x"12c2", x"12c5", 
    x"12c8", x"12cb", x"12ce", x"12d1", x"12d4", x"12d7", x"12db", x"12de", 
    x"12e1", x"12e4", x"12e7", x"12ea", x"12ed", x"12f0", x"12f3", x"12f7", 
    x"12fa", x"12fd", x"1300", x"1303", x"1306", x"1309", x"130c", x"130f", 
    x"1312", x"1316", x"1319", x"131c", x"131f", x"1322", x"1325", x"1328", 
    x"132b", x"132e", x"1332", x"1335", x"1338", x"133b", x"133e", x"1341", 
    x"1344", x"1347", x"134a", x"134d", x"1351", x"1354", x"1357", x"135a", 
    x"135d", x"1360", x"1363", x"1366", x"1369", x"136d", x"1370", x"1373", 
    x"1376", x"1379", x"137c", x"137f", x"1382", x"1385", x"1388", x"138c", 
    x"138f", x"1392", x"1395", x"1398", x"139b", x"139e", x"13a1", x"13a4", 
    x"13a8", x"13ab", x"13ae", x"13b1", x"13b4", x"13b7", x"13ba", x"13bd", 
    x"13c0", x"13c3", x"13c7", x"13ca", x"13cd", x"13d0", x"13d3", x"13d6", 
    x"13d9", x"13dc", x"13df", x"13e3", x"13e6", x"13e9", x"13ec", x"13ef", 
    x"13f2", x"13f5", x"13f8", x"13fb", x"13fe", x"1402", x"1405", x"1408", 
    x"140b", x"140e", x"1411", x"1414", x"1417", x"141a", x"141d", x"1421", 
    x"1424", x"1427", x"142a", x"142d", x"1430", x"1433", x"1436", x"1439", 
    x"143c", x"1440", x"1443", x"1446", x"1449", x"144c", x"144f", x"1452", 
    x"1455", x"1458", x"145c", x"145f", x"1462", x"1465", x"1468", x"146b", 
    x"146e", x"1471", x"1474", x"1477", x"147b", x"147e", x"1481", x"1484", 
    x"1487", x"148a", x"148d", x"1490", x"1493", x"1496", x"149a", x"149d", 
    x"14a0", x"14a3", x"14a6", x"14a9", x"14ac", x"14af", x"14b2", x"14b5", 
    x"14b9", x"14bc", x"14bf", x"14c2", x"14c5", x"14c8", x"14cb", x"14ce", 
    x"14d1", x"14d4", x"14d8", x"14db", x"14de", x"14e1", x"14e4", x"14e7", 
    x"14ea", x"14ed", x"14f0", x"14f3", x"14f7", x"14fa", x"14fd", x"1500", 
    x"1503", x"1506", x"1509", x"150c", x"150f", x"1512", x"1516", x"1519", 
    x"151c", x"151f", x"1522", x"1525", x"1528", x"152b", x"152e", x"1531", 
    x"1534", x"1538", x"153b", x"153e", x"1541", x"1544", x"1547", x"154a", 
    x"154d", x"1550", x"1553", x"1557", x"155a", x"155d", x"1560", x"1563", 
    x"1566", x"1569", x"156c", x"156f", x"1572", x"1576", x"1579", x"157c", 
    x"157f", x"1582", x"1585", x"1588", x"158b", x"158e", x"1591", x"1595", 
    x"1598", x"159b", x"159e", x"15a1", x"15a4", x"15a7", x"15aa", x"15ad", 
    x"15b0", x"15b3", x"15b7", x"15ba", x"15bd", x"15c0", x"15c3", x"15c6", 
    x"15c9", x"15cc", x"15cf", x"15d2", x"15d6", x"15d9", x"15dc", x"15df", 
    x"15e2", x"15e5", x"15e8", x"15eb", x"15ee", x"15f1", x"15f4", x"15f8", 
    x"15fb", x"15fe", x"1601", x"1604", x"1607", x"160a", x"160d", x"1610", 
    x"1613", x"1617", x"161a", x"161d", x"1620", x"1623", x"1626", x"1629", 
    x"162c", x"162f", x"1632", x"1635", x"1639", x"163c", x"163f", x"1642", 
    x"1645", x"1648", x"164b", x"164e", x"1651", x"1654", x"1657", x"165b", 
    x"165e", x"1661", x"1664", x"1667", x"166a", x"166d", x"1670", x"1673", 
    x"1676", x"167a", x"167d", x"1680", x"1683", x"1686", x"1689", x"168c", 
    x"168f", x"1692", x"1695", x"1698", x"169c", x"169f", x"16a2", x"16a5", 
    x"16a8", x"16ab", x"16ae", x"16b1", x"16b4", x"16b7", x"16ba", x"16be", 
    x"16c1", x"16c4", x"16c7", x"16ca", x"16cd", x"16d0", x"16d3", x"16d6", 
    x"16d9", x"16dc", x"16e0", x"16e3", x"16e6", x"16e9", x"16ec", x"16ef", 
    x"16f2", x"16f5", x"16f8", x"16fb", x"16fe", x"1702", x"1705", x"1708", 
    x"170b", x"170e", x"1711", x"1714", x"1717", x"171a", x"171d", x"1720", 
    x"1724", x"1727", x"172a", x"172d", x"1730", x"1733", x"1736", x"1739", 
    x"173c", x"173f", x"1742", x"1746", x"1749", x"174c", x"174f", x"1752", 
    x"1755", x"1758", x"175b", x"175e", x"1761", x"1764", x"1767", x"176b", 
    x"176e", x"1771", x"1774", x"1777", x"177a", x"177d", x"1780", x"1783", 
    x"1786", x"1789", x"178d", x"1790", x"1793", x"1796", x"1799", x"179c", 
    x"179f", x"17a2", x"17a5", x"17a8", x"17ab", x"17af", x"17b2", x"17b5", 
    x"17b8", x"17bb", x"17be", x"17c1", x"17c4", x"17c7", x"17ca", x"17cd", 
    x"17d0", x"17d4", x"17d7", x"17da", x"17dd", x"17e0", x"17e3", x"17e6", 
    x"17e9", x"17ec", x"17ef", x"17f2", x"17f6", x"17f9", x"17fc", x"17ff", 
    x"1802", x"1805", x"1808", x"180b", x"180e", x"1811", x"1814", x"1817", 
    x"181b", x"181e", x"1821", x"1824", x"1827", x"182a", x"182d", x"1830", 
    x"1833", x"1836", x"1839", x"183c", x"1840", x"1843", x"1846", x"1849", 
    x"184c", x"184f", x"1852", x"1855", x"1858", x"185b", x"185e", x"1861", 
    x"1865", x"1868", x"186b", x"186e", x"1871", x"1874", x"1877", x"187a", 
    x"187d", x"1880", x"1883", x"1886", x"188a", x"188d", x"1890", x"1893", 
    x"1896", x"1899", x"189c", x"189f", x"18a2", x"18a5", x"18a8", x"18ab", 
    x"18af", x"18b2", x"18b5", x"18b8", x"18bb", x"18be", x"18c1", x"18c4", 
    x"18c7", x"18ca", x"18cd", x"18d0", x"18d4", x"18d7", x"18da", x"18dd", 
    x"18e0", x"18e3", x"18e6", x"18e9", x"18ec", x"18ef", x"18f2", x"18f5", 
    x"18f9", x"18fc", x"18ff", x"1902", x"1905", x"1908", x"190b", x"190e", 
    x"1911", x"1914", x"1917", x"191a", x"191d", x"1921", x"1924", x"1927", 
    x"192a", x"192d", x"1930", x"1933", x"1936", x"1939", x"193c", x"193f", 
    x"1942", x"1946", x"1949", x"194c", x"194f", x"1952", x"1955", x"1958", 
    x"195b", x"195e", x"1961", x"1964", x"1967", x"196a", x"196e", x"1971", 
    x"1974", x"1977", x"197a", x"197d", x"1980", x"1983", x"1986", x"1989", 
    x"198c", x"198f", x"1993", x"1996", x"1999", x"199c", x"199f", x"19a2", 
    x"19a5", x"19a8", x"19ab", x"19ae", x"19b1", x"19b4", x"19b7", x"19bb", 
    x"19be", x"19c1", x"19c4", x"19c7", x"19ca", x"19cd", x"19d0", x"19d3", 
    x"19d6", x"19d9", x"19dc", x"19df", x"19e3", x"19e6", x"19e9", x"19ec", 
    x"19ef", x"19f2", x"19f5", x"19f8", x"19fb", x"19fe", x"1a01", x"1a04", 
    x"1a07", x"1a0b", x"1a0e", x"1a11", x"1a14", x"1a17", x"1a1a", x"1a1d", 
    x"1a20", x"1a23", x"1a26", x"1a29", x"1a2c", x"1a2f", x"1a32", x"1a36", 
    x"1a39", x"1a3c", x"1a3f", x"1a42", x"1a45", x"1a48", x"1a4b", x"1a4e", 
    x"1a51", x"1a54", x"1a57", x"1a5a", x"1a5e", x"1a61", x"1a64", x"1a67", 
    x"1a6a", x"1a6d", x"1a70", x"1a73", x"1a76", x"1a79", x"1a7c", x"1a7f", 
    x"1a82", x"1a85", x"1a89", x"1a8c", x"1a8f", x"1a92", x"1a95", x"1a98", 
    x"1a9b", x"1a9e", x"1aa1", x"1aa4", x"1aa7", x"1aaa", x"1aad", x"1ab1", 
    x"1ab4", x"1ab7", x"1aba", x"1abd", x"1ac0", x"1ac3", x"1ac6", x"1ac9", 
    x"1acc", x"1acf", x"1ad2", x"1ad5", x"1ad8", x"1adc", x"1adf", x"1ae2", 
    x"1ae5", x"1ae8", x"1aeb", x"1aee", x"1af1", x"1af4", x"1af7", x"1afa", 
    x"1afd", x"1b00", x"1b03", x"1b07", x"1b0a", x"1b0d", x"1b10", x"1b13", 
    x"1b16", x"1b19", x"1b1c", x"1b1f", x"1b22", x"1b25", x"1b28", x"1b2b", 
    x"1b2e", x"1b31", x"1b35", x"1b38", x"1b3b", x"1b3e", x"1b41", x"1b44", 
    x"1b47", x"1b4a", x"1b4d", x"1b50", x"1b53", x"1b56", x"1b59", x"1b5c", 
    x"1b60", x"1b63", x"1b66", x"1b69", x"1b6c", x"1b6f", x"1b72", x"1b75", 
    x"1b78", x"1b7b", x"1b7e", x"1b81", x"1b84", x"1b87", x"1b8a", x"1b8e", 
    x"1b91", x"1b94", x"1b97", x"1b9a", x"1b9d", x"1ba0", x"1ba3", x"1ba6", 
    x"1ba9", x"1bac", x"1baf", x"1bb2", x"1bb5", x"1bb9", x"1bbc", x"1bbf", 
    x"1bc2", x"1bc5", x"1bc8", x"1bcb", x"1bce", x"1bd1", x"1bd4", x"1bd7", 
    x"1bda", x"1bdd", x"1be0", x"1be3", x"1be7", x"1bea", x"1bed", x"1bf0", 
    x"1bf3", x"1bf6", x"1bf9", x"1bfc", x"1bff", x"1c02", x"1c05", x"1c08", 
    x"1c0b", x"1c0e", x"1c11", x"1c14", x"1c18", x"1c1b", x"1c1e", x"1c21", 
    x"1c24", x"1c27", x"1c2a", x"1c2d", x"1c30", x"1c33", x"1c36", x"1c39", 
    x"1c3c", x"1c3f", x"1c42", x"1c46", x"1c49", x"1c4c", x"1c4f", x"1c52", 
    x"1c55", x"1c58", x"1c5b", x"1c5e", x"1c61", x"1c64", x"1c67", x"1c6a", 
    x"1c6d", x"1c70", x"1c73", x"1c77", x"1c7a", x"1c7d", x"1c80", x"1c83", 
    x"1c86", x"1c89", x"1c8c", x"1c8f", x"1c92", x"1c95", x"1c98", x"1c9b", 
    x"1c9e", x"1ca1", x"1ca4", x"1ca8", x"1cab", x"1cae", x"1cb1", x"1cb4", 
    x"1cb7", x"1cba", x"1cbd", x"1cc0", x"1cc3", x"1cc6", x"1cc9", x"1ccc", 
    x"1ccf", x"1cd2", x"1cd5", x"1cd9", x"1cdc", x"1cdf", x"1ce2", x"1ce5", 
    x"1ce8", x"1ceb", x"1cee", x"1cf1", x"1cf4", x"1cf7", x"1cfa", x"1cfd", 
    x"1d00", x"1d03", x"1d06", x"1d09", x"1d0d", x"1d10", x"1d13", x"1d16", 
    x"1d19", x"1d1c", x"1d1f", x"1d22", x"1d25", x"1d28", x"1d2b", x"1d2e", 
    x"1d31", x"1d34", x"1d37", x"1d3a", x"1d3d", x"1d41", x"1d44", x"1d47", 
    x"1d4a", x"1d4d", x"1d50", x"1d53", x"1d56", x"1d59", x"1d5c", x"1d5f", 
    x"1d62", x"1d65", x"1d68", x"1d6b", x"1d6e", x"1d71", x"1d75", x"1d78", 
    x"1d7b", x"1d7e", x"1d81", x"1d84", x"1d87", x"1d8a", x"1d8d", x"1d90", 
    x"1d93", x"1d96", x"1d99", x"1d9c", x"1d9f", x"1da2", x"1da5", x"1da8", 
    x"1dac", x"1daf", x"1db2", x"1db5", x"1db8", x"1dbb", x"1dbe", x"1dc1", 
    x"1dc4", x"1dc7", x"1dca", x"1dcd", x"1dd0", x"1dd3", x"1dd6", x"1dd9", 
    x"1ddc", x"1ddf", x"1de3", x"1de6", x"1de9", x"1dec", x"1def", x"1df2", 
    x"1df5", x"1df8", x"1dfb", x"1dfe", x"1e01", x"1e04", x"1e07", x"1e0a", 
    x"1e0d", x"1e10", x"1e13", x"1e16", x"1e19", x"1e1d", x"1e20", x"1e23", 
    x"1e26", x"1e29", x"1e2c", x"1e2f", x"1e32", x"1e35", x"1e38", x"1e3b", 
    x"1e3e", x"1e41", x"1e44", x"1e47", x"1e4a", x"1e4d", x"1e50", x"1e54", 
    x"1e57", x"1e5a", x"1e5d", x"1e60", x"1e63", x"1e66", x"1e69", x"1e6c", 
    x"1e6f", x"1e72", x"1e75", x"1e78", x"1e7b", x"1e7e", x"1e81", x"1e84", 
    x"1e87", x"1e8a", x"1e8d", x"1e91", x"1e94", x"1e97", x"1e9a", x"1e9d", 
    x"1ea0", x"1ea3", x"1ea6", x"1ea9", x"1eac", x"1eaf", x"1eb2", x"1eb5", 
    x"1eb8", x"1ebb", x"1ebe", x"1ec1", x"1ec4", x"1ec7", x"1eca", x"1ece", 
    x"1ed1", x"1ed4", x"1ed7", x"1eda", x"1edd", x"1ee0", x"1ee3", x"1ee6", 
    x"1ee9", x"1eec", x"1eef", x"1ef2", x"1ef5", x"1ef8", x"1efb", x"1efe", 
    x"1f01", x"1f04", x"1f07", x"1f0a", x"1f0e", x"1f11", x"1f14", x"1f17", 
    x"1f1a", x"1f1d", x"1f20", x"1f23", x"1f26", x"1f29", x"1f2c", x"1f2f", 
    x"1f32", x"1f35", x"1f38", x"1f3b", x"1f3e", x"1f41", x"1f44", x"1f47", 
    x"1f4a", x"1f4e", x"1f51", x"1f54", x"1f57", x"1f5a", x"1f5d", x"1f60", 
    x"1f63", x"1f66", x"1f69", x"1f6c", x"1f6f", x"1f72", x"1f75", x"1f78", 
    x"1f7b", x"1f7e", x"1f81", x"1f84", x"1f87", x"1f8a", x"1f8d", x"1f91", 
    x"1f94", x"1f97", x"1f9a", x"1f9d", x"1fa0", x"1fa3", x"1fa6", x"1fa9", 
    x"1fac", x"1faf", x"1fb2", x"1fb5", x"1fb8", x"1fbb", x"1fbe", x"1fc1", 
    x"1fc4", x"1fc7", x"1fca", x"1fcd", x"1fd0", x"1fd3", x"1fd7", x"1fda", 
    x"1fdd", x"1fe0", x"1fe3", x"1fe6", x"1fe9", x"1fec", x"1fef", x"1ff2", 
    x"1ff5", x"1ff8", x"1ffb", x"1ffe", x"2001", x"2004", x"2007", x"200a", 
    x"200d", x"2010", x"2013", x"2016", x"2019", x"201c", x"2020", x"2023", 
    x"2026", x"2029", x"202c", x"202f", x"2032", x"2035", x"2038", x"203b", 
    x"203e", x"2041", x"2044", x"2047", x"204a", x"204d", x"2050", x"2053", 
    x"2056", x"2059", x"205c", x"205f", x"2062", x"2065", x"2068", x"206c", 
    x"206f", x"2072", x"2075", x"2078", x"207b", x"207e", x"2081", x"2084", 
    x"2087", x"208a", x"208d", x"2090", x"2093", x"2096", x"2099", x"209c", 
    x"209f", x"20a2", x"20a5", x"20a8", x"20ab", x"20ae", x"20b1", x"20b4", 
    x"20b7", x"20bb", x"20be", x"20c1", x"20c4", x"20c7", x"20ca", x"20cd", 
    x"20d0", x"20d3", x"20d6", x"20d9", x"20dc", x"20df", x"20e2", x"20e5", 
    x"20e8", x"20eb", x"20ee", x"20f1", x"20f4", x"20f7", x"20fa", x"20fd", 
    x"2100", x"2103", x"2106", x"2109", x"210c", x"2110", x"2113", x"2116", 
    x"2119", x"211c", x"211f", x"2122", x"2125", x"2128", x"212b", x"212e", 
    x"2131", x"2134", x"2137", x"213a", x"213d", x"2140", x"2143", x"2146", 
    x"2149", x"214c", x"214f", x"2152", x"2155", x"2158", x"215b", x"215e", 
    x"2161", x"2164", x"2168", x"216b", x"216e", x"2171", x"2174", x"2177", 
    x"217a", x"217d", x"2180", x"2183", x"2186", x"2189", x"218c", x"218f", 
    x"2192", x"2195", x"2198", x"219b", x"219e", x"21a1", x"21a4", x"21a7", 
    x"21aa", x"21ad", x"21b0", x"21b3", x"21b6", x"21b9", x"21bc", x"21bf", 
    x"21c2", x"21c5", x"21c9", x"21cc", x"21cf", x"21d2", x"21d5", x"21d8", 
    x"21db", x"21de", x"21e1", x"21e4", x"21e7", x"21ea", x"21ed", x"21f0", 
    x"21f3", x"21f6", x"21f9", x"21fc", x"21ff", x"2202", x"2205", x"2208", 
    x"220b", x"220e", x"2211", x"2214", x"2217", x"221a", x"221d", x"2220", 
    x"2223", x"2226", x"2229", x"222c", x"222f", x"2233", x"2236", x"2239", 
    x"223c", x"223f", x"2242", x"2245", x"2248", x"224b", x"224e", x"2251", 
    x"2254", x"2257", x"225a", x"225d", x"2260", x"2263", x"2266", x"2269", 
    x"226c", x"226f", x"2272", x"2275", x"2278", x"227b", x"227e", x"2281", 
    x"2284", x"2287", x"228a", x"228d", x"2290", x"2293", x"2296", x"2299", 
    x"229c", x"229f", x"22a2", x"22a5", x"22a9", x"22ac", x"22af", x"22b2", 
    x"22b5", x"22b8", x"22bb", x"22be", x"22c1", x"22c4", x"22c7", x"22ca", 
    x"22cd", x"22d0", x"22d3", x"22d6", x"22d9", x"22dc", x"22df", x"22e2", 
    x"22e5", x"22e8", x"22eb", x"22ee", x"22f1", x"22f4", x"22f7", x"22fa", 
    x"22fd", x"2300", x"2303", x"2306", x"2309", x"230c", x"230f", x"2312", 
    x"2315", x"2318", x"231b", x"231e", x"2321", x"2324", x"2327", x"232a", 
    x"232e", x"2331", x"2334", x"2337", x"233a", x"233d", x"2340", x"2343", 
    x"2346", x"2349", x"234c", x"234f", x"2352", x"2355", x"2358", x"235b", 
    x"235e", x"2361", x"2364", x"2367", x"236a", x"236d", x"2370", x"2373", 
    x"2376", x"2379", x"237c", x"237f", x"2382", x"2385", x"2388", x"238b", 
    x"238e", x"2391", x"2394", x"2397", x"239a", x"239d", x"23a0", x"23a3", 
    x"23a6", x"23a9", x"23ac", x"23af", x"23b2", x"23b5", x"23b8", x"23bb", 
    x"23be", x"23c1", x"23c4", x"23c7", x"23ca", x"23cd", x"23d0", x"23d4", 
    x"23d7", x"23da", x"23dd", x"23e0", x"23e3", x"23e6", x"23e9", x"23ec", 
    x"23ef", x"23f2", x"23f5", x"23f8", x"23fb", x"23fe", x"2401", x"2404", 
    x"2407", x"240a", x"240d", x"2410", x"2413", x"2416", x"2419", x"241c", 
    x"241f", x"2422", x"2425", x"2428", x"242b", x"242e", x"2431", x"2434", 
    x"2437", x"243a", x"243d", x"2440", x"2443", x"2446", x"2449", x"244c", 
    x"244f", x"2452", x"2455", x"2458", x"245b", x"245e", x"2461", x"2464", 
    x"2467", x"246a", x"246d", x"2470", x"2473", x"2476", x"2479", x"247c", 
    x"247f", x"2482", x"2485", x"2488", x"248b", x"248e", x"2491", x"2494", 
    x"2497", x"249a", x"249d", x"24a0", x"24a3", x"24a6", x"24a9", x"24ac", 
    x"24af", x"24b2", x"24b5", x"24b8", x"24bb", x"24be", x"24c1", x"24c5", 
    x"24c8", x"24cb", x"24ce", x"24d1", x"24d4", x"24d7", x"24da", x"24dd", 
    x"24e0", x"24e3", x"24e6", x"24e9", x"24ec", x"24ef", x"24f2", x"24f5", 
    x"24f8", x"24fb", x"24fe", x"2501", x"2504", x"2507", x"250a", x"250d", 
    x"2510", x"2513", x"2516", x"2519", x"251c", x"251f", x"2522", x"2525", 
    x"2528", x"252b", x"252e", x"2531", x"2534", x"2537", x"253a", x"253d", 
    x"2540", x"2543", x"2546", x"2549", x"254c", x"254f", x"2552", x"2555", 
    x"2558", x"255b", x"255e", x"2561", x"2564", x"2567", x"256a", x"256d", 
    x"2570", x"2573", x"2576", x"2579", x"257c", x"257f", x"2582", x"2585", 
    x"2588", x"258b", x"258e", x"2591", x"2594", x"2597", x"259a", x"259d", 
    x"25a0", x"25a3", x"25a6", x"25a9", x"25ac", x"25af", x"25b2", x"25b5", 
    x"25b8", x"25bb", x"25be", x"25c1", x"25c4", x"25c7", x"25ca", x"25cd", 
    x"25d0", x"25d3", x"25d6", x"25d9", x"25dc", x"25df", x"25e2", x"25e5", 
    x"25e8", x"25eb", x"25ee", x"25f1", x"25f4", x"25f7", x"25fa", x"25fd", 
    x"2600", x"2603", x"2606", x"2609", x"260c", x"260f", x"2612", x"2615", 
    x"2618", x"261b", x"261e", x"2621", x"2624", x"2627", x"262a", x"262d", 
    x"2630", x"2633", x"2636", x"2639", x"263c", x"263f", x"2642", x"2645", 
    x"2648", x"264b", x"264e", x"2651", x"2654", x"2657", x"265a", x"265d", 
    x"2660", x"2663", x"2666", x"2669", x"266c", x"266f", x"2672", x"2675", 
    x"2678", x"267b", x"267e", x"2681", x"2684", x"2687", x"268a", x"268d", 
    x"2690", x"2693", x"2696", x"2699", x"269c", x"269f", x"26a2", x"26a5", 
    x"26a8", x"26ab", x"26ae", x"26b1", x"26b4", x"26b7", x"26ba", x"26bd", 
    x"26c0", x"26c3", x"26c6", x"26c9", x"26cc", x"26cf", x"26d2", x"26d5", 
    x"26d8", x"26db", x"26de", x"26e1", x"26e4", x"26e7", x"26ea", x"26ed", 
    x"26f0", x"26f3", x"26f6", x"26f9", x"26fc", x"26ff", x"2702", x"2705", 
    x"2708", x"270b", x"270e", x"2711", x"2714", x"2717", x"271a", x"271d", 
    x"2720", x"2723", x"2726", x"2729", x"272c", x"272f", x"2731", x"2734", 
    x"2737", x"273a", x"273d", x"2740", x"2743", x"2746", x"2749", x"274c", 
    x"274f", x"2752", x"2755", x"2758", x"275b", x"275e", x"2761", x"2764", 
    x"2767", x"276a", x"276d", x"2770", x"2773", x"2776", x"2779", x"277c", 
    x"277f", x"2782", x"2785", x"2788", x"278b", x"278e", x"2791", x"2794", 
    x"2797", x"279a", x"279d", x"27a0", x"27a3", x"27a6", x"27a9", x"27ac", 
    x"27af", x"27b2", x"27b5", x"27b8", x"27bb", x"27be", x"27c1", x"27c4", 
    x"27c7", x"27ca", x"27cd", x"27d0", x"27d3", x"27d6", x"27d9", x"27dc", 
    x"27df", x"27e2", x"27e5", x"27e8", x"27eb", x"27ee", x"27f1", x"27f4", 
    x"27f7", x"27fa", x"27fd", x"2800", x"2803", x"2806", x"2809", x"280c", 
    x"280f", x"2812", x"2815", x"2817", x"281a", x"281d", x"2820", x"2823", 
    x"2826", x"2829", x"282c", x"282f", x"2832", x"2835", x"2838", x"283b", 
    x"283e", x"2841", x"2844", x"2847", x"284a", x"284d", x"2850", x"2853", 
    x"2856", x"2859", x"285c", x"285f", x"2862", x"2865", x"2868", x"286b", 
    x"286e", x"2871", x"2874", x"2877", x"287a", x"287d", x"2880", x"2883", 
    x"2886", x"2889", x"288c", x"288f", x"2892", x"2895", x"2898", x"289b", 
    x"289e", x"28a1", x"28a4", x"28a7", x"28aa", x"28ad", x"28b0", x"28b3", 
    x"28b5", x"28b8", x"28bb", x"28be", x"28c1", x"28c4", x"28c7", x"28ca", 
    x"28cd", x"28d0", x"28d3", x"28d6", x"28d9", x"28dc", x"28df", x"28e2", 
    x"28e5", x"28e8", x"28eb", x"28ee", x"28f1", x"28f4", x"28f7", x"28fa", 
    x"28fd", x"2900", x"2903", x"2906", x"2909", x"290c", x"290f", x"2912", 
    x"2915", x"2918", x"291b", x"291e", x"2921", x"2924", x"2927", x"292a", 
    x"292d", x"2930", x"2932", x"2935", x"2938", x"293b", x"293e", x"2941", 
    x"2944", x"2947", x"294a", x"294d", x"2950", x"2953", x"2956", x"2959", 
    x"295c", x"295f", x"2962", x"2965", x"2968", x"296b", x"296e", x"2971", 
    x"2974", x"2977", x"297a", x"297d", x"2980", x"2983", x"2986", x"2989", 
    x"298c", x"298f", x"2992", x"2995", x"2998", x"299b", x"299e", x"29a0", 
    x"29a3", x"29a6", x"29a9", x"29ac", x"29af", x"29b2", x"29b5", x"29b8", 
    x"29bb", x"29be", x"29c1", x"29c4", x"29c7", x"29ca", x"29cd", x"29d0", 
    x"29d3", x"29d6", x"29d9", x"29dc", x"29df", x"29e2", x"29e5", x"29e8", 
    x"29eb", x"29ee", x"29f1", x"29f4", x"29f7", x"29fa", x"29fd", x"29ff", 
    x"2a02", x"2a05", x"2a08", x"2a0b", x"2a0e", x"2a11", x"2a14", x"2a17", 
    x"2a1a", x"2a1d", x"2a20", x"2a23", x"2a26", x"2a29", x"2a2c", x"2a2f", 
    x"2a32", x"2a35", x"2a38", x"2a3b", x"2a3e", x"2a41", x"2a44", x"2a47", 
    x"2a4a", x"2a4d", x"2a50", x"2a53", x"2a56", x"2a58", x"2a5b", x"2a5e", 
    x"2a61", x"2a64", x"2a67", x"2a6a", x"2a6d", x"2a70", x"2a73", x"2a76", 
    x"2a79", x"2a7c", x"2a7f", x"2a82", x"2a85", x"2a88", x"2a8b", x"2a8e", 
    x"2a91", x"2a94", x"2a97", x"2a9a", x"2a9d", x"2aa0", x"2aa3", x"2aa6", 
    x"2aa8", x"2aab", x"2aae", x"2ab1", x"2ab4", x"2ab7", x"2aba", x"2abd", 
    x"2ac0", x"2ac3", x"2ac6", x"2ac9", x"2acc", x"2acf", x"2ad2", x"2ad5", 
    x"2ad8", x"2adb", x"2ade", x"2ae1", x"2ae4", x"2ae7", x"2aea", x"2aed", 
    x"2af0", x"2af2", x"2af5", x"2af8", x"2afb", x"2afe", x"2b01", x"2b04", 
    x"2b07", x"2b0a", x"2b0d", x"2b10", x"2b13", x"2b16", x"2b19", x"2b1c", 
    x"2b1f", x"2b22", x"2b25", x"2b28", x"2b2b", x"2b2e", x"2b31", x"2b34", 
    x"2b37", x"2b39", x"2b3c", x"2b3f", x"2b42", x"2b45", x"2b48", x"2b4b", 
    x"2b4e", x"2b51", x"2b54", x"2b57", x"2b5a", x"2b5d", x"2b60", x"2b63", 
    x"2b66", x"2b69", x"2b6c", x"2b6f", x"2b72", x"2b75", x"2b78", x"2b7b", 
    x"2b7d", x"2b80", x"2b83", x"2b86", x"2b89", x"2b8c", x"2b8f", x"2b92", 
    x"2b95", x"2b98", x"2b9b", x"2b9e", x"2ba1", x"2ba4", x"2ba7", x"2baa", 
    x"2bad", x"2bb0", x"2bb3", x"2bb6", x"2bb9", x"2bbb", x"2bbe", x"2bc1", 
    x"2bc4", x"2bc7", x"2bca", x"2bcd", x"2bd0", x"2bd3", x"2bd6", x"2bd9", 
    x"2bdc", x"2bdf", x"2be2", x"2be5", x"2be8", x"2beb", x"2bee", x"2bf1", 
    x"2bf4", x"2bf7", x"2bf9", x"2bfc", x"2bff", x"2c02", x"2c05", x"2c08", 
    x"2c0b", x"2c0e", x"2c11", x"2c14", x"2c17", x"2c1a", x"2c1d", x"2c20", 
    x"2c23", x"2c26", x"2c29", x"2c2c", x"2c2f", x"2c32", x"2c34", x"2c37", 
    x"2c3a", x"2c3d", x"2c40", x"2c43", x"2c46", x"2c49", x"2c4c", x"2c4f", 
    x"2c52", x"2c55", x"2c58", x"2c5b", x"2c5e", x"2c61", x"2c64", x"2c67", 
    x"2c6a", x"2c6c", x"2c6f", x"2c72", x"2c75", x"2c78", x"2c7b", x"2c7e", 
    x"2c81", x"2c84", x"2c87", x"2c8a", x"2c8d", x"2c90", x"2c93", x"2c96", 
    x"2c99", x"2c9c", x"2c9f", x"2ca1", x"2ca4", x"2ca7", x"2caa", x"2cad", 
    x"2cb0", x"2cb3", x"2cb6", x"2cb9", x"2cbc", x"2cbf", x"2cc2", x"2cc5", 
    x"2cc8", x"2ccb", x"2cce", x"2cd1", x"2cd4", x"2cd6", x"2cd9", x"2cdc", 
    x"2cdf", x"2ce2", x"2ce5", x"2ce8", x"2ceb", x"2cee", x"2cf1", x"2cf4", 
    x"2cf7", x"2cfa", x"2cfd", x"2d00", x"2d03", x"2d06", x"2d08", x"2d0b", 
    x"2d0e", x"2d11", x"2d14", x"2d17", x"2d1a", x"2d1d", x"2d20", x"2d23", 
    x"2d26", x"2d29", x"2d2c", x"2d2f", x"2d32", x"2d35", x"2d37", x"2d3a", 
    x"2d3d", x"2d40", x"2d43", x"2d46", x"2d49", x"2d4c", x"2d4f", x"2d52", 
    x"2d55", x"2d58", x"2d5b", x"2d5e", x"2d61", x"2d64", x"2d67", x"2d69", 
    x"2d6c", x"2d6f", x"2d72", x"2d75", x"2d78", x"2d7b", x"2d7e", x"2d81", 
    x"2d84", x"2d87", x"2d8a", x"2d8d", x"2d90", x"2d93", x"2d95", x"2d98", 
    x"2d9b", x"2d9e", x"2da1", x"2da4", x"2da7", x"2daa", x"2dad", x"2db0", 
    x"2db3", x"2db6", x"2db9", x"2dbc", x"2dbf", x"2dc2", x"2dc4", x"2dc7", 
    x"2dca", x"2dcd", x"2dd0", x"2dd3", x"2dd6", x"2dd9", x"2ddc", x"2ddf", 
    x"2de2", x"2de5", x"2de8", x"2deb", x"2dee", x"2df0", x"2df3", x"2df6", 
    x"2df9", x"2dfc", x"2dff", x"2e02", x"2e05", x"2e08", x"2e0b", x"2e0e", 
    x"2e11", x"2e14", x"2e17", x"2e19", x"2e1c", x"2e1f", x"2e22", x"2e25", 
    x"2e28", x"2e2b", x"2e2e", x"2e31", x"2e34", x"2e37", x"2e3a", x"2e3d", 
    x"2e40", x"2e42", x"2e45", x"2e48", x"2e4b", x"2e4e", x"2e51", x"2e54", 
    x"2e57", x"2e5a", x"2e5d", x"2e60", x"2e63", x"2e66", x"2e69", x"2e6b", 
    x"2e6e", x"2e71", x"2e74", x"2e77", x"2e7a", x"2e7d", x"2e80", x"2e83", 
    x"2e86", x"2e89", x"2e8c", x"2e8f", x"2e92", x"2e94", x"2e97", x"2e9a", 
    x"2e9d", x"2ea0", x"2ea3", x"2ea6", x"2ea9", x"2eac", x"2eaf", x"2eb2", 
    x"2eb5", x"2eb8", x"2eba", x"2ebd", x"2ec0", x"2ec3", x"2ec6", x"2ec9", 
    x"2ecc", x"2ecf", x"2ed2", x"2ed5", x"2ed8", x"2edb", x"2ede", x"2ee1", 
    x"2ee3", x"2ee6", x"2ee9", x"2eec", x"2eef", x"2ef2", x"2ef5", x"2ef8", 
    x"2efb", x"2efe", x"2f01", x"2f04", x"2f06", x"2f09", x"2f0c", x"2f0f", 
    x"2f12", x"2f15", x"2f18", x"2f1b", x"2f1e", x"2f21", x"2f24", x"2f27", 
    x"2f2a", x"2f2c", x"2f2f", x"2f32", x"2f35", x"2f38", x"2f3b", x"2f3e", 
    x"2f41", x"2f44", x"2f47", x"2f4a", x"2f4d", x"2f50", x"2f52", x"2f55", 
    x"2f58", x"2f5b", x"2f5e", x"2f61", x"2f64", x"2f67", x"2f6a", x"2f6d", 
    x"2f70", x"2f73", x"2f75", x"2f78", x"2f7b", x"2f7e", x"2f81", x"2f84", 
    x"2f87", x"2f8a", x"2f8d", x"2f90", x"2f93", x"2f96", x"2f98", x"2f9b", 
    x"2f9e", x"2fa1", x"2fa4", x"2fa7", x"2faa", x"2fad", x"2fb0", x"2fb3", 
    x"2fb6", x"2fb9", x"2fbb", x"2fbe", x"2fc1", x"2fc4", x"2fc7", x"2fca", 
    x"2fcd", x"2fd0", x"2fd3", x"2fd6", x"2fd9", x"2fdb", x"2fde", x"2fe1", 
    x"2fe4", x"2fe7", x"2fea", x"2fed", x"2ff0", x"2ff3", x"2ff6", x"2ff9", 
    x"2ffc", x"2ffe", x"3001", x"3004", x"3007", x"300a", x"300d", x"3010", 
    x"3013", x"3016", x"3019", x"301c", x"301e", x"3021", x"3024", x"3027", 
    x"302a", x"302d", x"3030", x"3033", x"3036", x"3039", x"303c", x"303e", 
    x"3041", x"3044", x"3047", x"304a", x"304d", x"3050", x"3053", x"3056", 
    x"3059", x"305c", x"305e", x"3061", x"3064", x"3067", x"306a", x"306d", 
    x"3070", x"3073", x"3076", x"3079", x"307c", x"307e", x"3081", x"3084", 
    x"3087", x"308a", x"308d", x"3090", x"3093", x"3096", x"3099", x"309c", 
    x"309e", x"30a1", x"30a4", x"30a7", x"30aa", x"30ad", x"30b0", x"30b3", 
    x"30b6", x"30b9", x"30bc", x"30be", x"30c1", x"30c4", x"30c7", x"30ca", 
    x"30cd", x"30d0", x"30d3", x"30d6", x"30d9", x"30db", x"30de", x"30e1", 
    x"30e4", x"30e7", x"30ea", x"30ed", x"30f0", x"30f3", x"30f6", x"30f8", 
    x"30fb", x"30fe", x"3101", x"3104", x"3107", x"310a", x"310d", x"3110", 
    x"3113", x"3116", x"3118", x"311b", x"311e", x"3121", x"3124", x"3127", 
    x"312a", x"312d", x"3130", x"3133", x"3135", x"3138", x"313b", x"313e", 
    x"3141", x"3144", x"3147", x"314a", x"314d", x"3150", x"3152", x"3155", 
    x"3158", x"315b", x"315e", x"3161", x"3164", x"3167", x"316a", x"316c", 
    x"316f", x"3172", x"3175", x"3178", x"317b", x"317e", x"3181", x"3184", 
    x"3187", x"3189", x"318c", x"318f", x"3192", x"3195", x"3198", x"319b", 
    x"319e", x"31a1", x"31a4", x"31a6", x"31a9", x"31ac", x"31af", x"31b2", 
    x"31b5", x"31b8", x"31bb", x"31be", x"31c0", x"31c3", x"31c6", x"31c9", 
    x"31cc", x"31cf", x"31d2", x"31d5", x"31d8", x"31db", x"31dd", x"31e0", 
    x"31e3", x"31e6", x"31e9", x"31ec", x"31ef", x"31f2", x"31f5", x"31f7", 
    x"31fa", x"31fd", x"3200", x"3203", x"3206", x"3209", x"320c", x"320f", 
    x"3211", x"3214", x"3217", x"321a", x"321d", x"3220", x"3223", x"3226", 
    x"3229", x"322b", x"322e", x"3231", x"3234", x"3237", x"323a", x"323d", 
    x"3240", x"3243", x"3246", x"3248", x"324b", x"324e", x"3251", x"3254", 
    x"3257", x"325a", x"325d", x"325f", x"3262", x"3265", x"3268", x"326b", 
    x"326e", x"3271", x"3274", x"3277", x"3279", x"327c", x"327f", x"3282", 
    x"3285", x"3288", x"328b", x"328e", x"3291", x"3293", x"3296", x"3299", 
    x"329c", x"329f", x"32a2", x"32a5", x"32a8", x"32ab", x"32ad", x"32b0", 
    x"32b3", x"32b6", x"32b9", x"32bc", x"32bf", x"32c2", x"32c5", x"32c7", 
    x"32ca", x"32cd", x"32d0", x"32d3", x"32d6", x"32d9", x"32dc", x"32de", 
    x"32e1", x"32e4", x"32e7", x"32ea", x"32ed", x"32f0", x"32f3", x"32f6", 
    x"32f8", x"32fb", x"32fe", x"3301", x"3304", x"3307", x"330a", x"330d", 
    x"330f", x"3312", x"3315", x"3318", x"331b", x"331e", x"3321", x"3324", 
    x"3326", x"3329", x"332c", x"332f", x"3332", x"3335", x"3338", x"333b", 
    x"333e", x"3340", x"3343", x"3346", x"3349", x"334c", x"334f", x"3352", 
    x"3355", x"3357", x"335a", x"335d", x"3360", x"3363", x"3366", x"3369", 
    x"336c", x"336e", x"3371", x"3374", x"3377", x"337a", x"337d", x"3380", 
    x"3383", x"3385", x"3388", x"338b", x"338e", x"3391", x"3394", x"3397", 
    x"339a", x"339c", x"339f", x"33a2", x"33a5", x"33a8", x"33ab", x"33ae", 
    x"33b1", x"33b3", x"33b6", x"33b9", x"33bc", x"33bf", x"33c2", x"33c5", 
    x"33c8", x"33ca", x"33cd", x"33d0", x"33d3", x"33d6", x"33d9", x"33dc", 
    x"33df", x"33e1", x"33e4", x"33e7", x"33ea", x"33ed", x"33f0", x"33f3", 
    x"33f6", x"33f8", x"33fb", x"33fe", x"3401", x"3404", x"3407", x"340a", 
    x"340c", x"340f", x"3412", x"3415", x"3418", x"341b", x"341e", x"3421", 
    x"3423", x"3426", x"3429", x"342c", x"342f", x"3432", x"3435", x"3438", 
    x"343a", x"343d", x"3440", x"3443", x"3446", x"3449", x"344c", x"344e", 
    x"3451", x"3454", x"3457", x"345a", x"345d", x"3460", x"3463", x"3465", 
    x"3468", x"346b", x"346e", x"3471", x"3474", x"3477", x"3479", x"347c", 
    x"347f", x"3482", x"3485", x"3488", x"348b", x"348e", x"3490", x"3493", 
    x"3496", x"3499", x"349c", x"349f", x"34a2", x"34a4", x"34a7", x"34aa", 
    x"34ad", x"34b0", x"34b3", x"34b6", x"34b8", x"34bb", x"34be", x"34c1", 
    x"34c4", x"34c7", x"34ca", x"34cc", x"34cf", x"34d2", x"34d5", x"34d8", 
    x"34db", x"34de", x"34e1", x"34e3", x"34e6", x"34e9", x"34ec", x"34ef", 
    x"34f2", x"34f5", x"34f7", x"34fa", x"34fd", x"3500", x"3503", x"3506", 
    x"3509", x"350b", x"350e", x"3511", x"3514", x"3517", x"351a", x"351d", 
    x"351f", x"3522", x"3525", x"3528", x"352b", x"352e", x"3531", x"3533", 
    x"3536", x"3539", x"353c", x"353f", x"3542", x"3545", x"3547", x"354a", 
    x"354d", x"3550", x"3553", x"3556", x"3559", x"355b", x"355e", x"3561", 
    x"3564", x"3567", x"356a", x"356d", x"356f", x"3572", x"3575", x"3578", 
    x"357b", x"357e", x"3581", x"3583", x"3586", x"3589", x"358c", x"358f", 
    x"3592", x"3595", x"3597", x"359a", x"359d", x"35a0", x"35a3", x"35a6", 
    x"35a8", x"35ab", x"35ae", x"35b1", x"35b4", x"35b7", x"35ba", x"35bc", 
    x"35bf", x"35c2", x"35c5", x"35c8", x"35cb", x"35ce", x"35d0", x"35d3", 
    x"35d6", x"35d9", x"35dc", x"35df", x"35e1", x"35e4", x"35e7", x"35ea", 
    x"35ed", x"35f0", x"35f3", x"35f5", x"35f8", x"35fb", x"35fe", x"3601", 
    x"3604", x"3607", x"3609", x"360c", x"360f", x"3612", x"3615", x"3618", 
    x"361a", x"361d", x"3620", x"3623", x"3626", x"3629", x"362c", x"362e", 
    x"3631", x"3634", x"3637", x"363a", x"363d", x"363f", x"3642", x"3645", 
    x"3648", x"364b", x"364e", x"3651", x"3653", x"3656", x"3659", x"365c", 
    x"365f", x"3662", x"3664", x"3667", x"366a", x"366d", x"3670", x"3673", 
    x"3676", x"3678", x"367b", x"367e", x"3681", x"3684", x"3687", x"3689", 
    x"368c", x"368f", x"3692", x"3695", x"3698", x"369a", x"369d", x"36a0", 
    x"36a3", x"36a6", x"36a9", x"36ab", x"36ae", x"36b1", x"36b4", x"36b7", 
    x"36ba", x"36bd", x"36bf", x"36c2", x"36c5", x"36c8", x"36cb", x"36ce", 
    x"36d0", x"36d3", x"36d6", x"36d9", x"36dc", x"36df", x"36e1", x"36e4", 
    x"36e7", x"36ea", x"36ed", x"36f0", x"36f2", x"36f5", x"36f8", x"36fb", 
    x"36fe", x"3701", x"3703", x"3706", x"3709", x"370c", x"370f", x"3712", 
    x"3715", x"3717", x"371a", x"371d", x"3720", x"3723", x"3726", x"3728", 
    x"372b", x"372e", x"3731", x"3734", x"3737", x"3739", x"373c", x"373f", 
    x"3742", x"3745", x"3748", x"374a", x"374d", x"3750", x"3753", x"3756", 
    x"3759", x"375b", x"375e", x"3761", x"3764", x"3767", x"376a", x"376c", 
    x"376f", x"3772", x"3775", x"3778", x"377b", x"377d", x"3780", x"3783", 
    x"3786", x"3789", x"378b", x"378e", x"3791", x"3794", x"3797", x"379a", 
    x"379c", x"379f", x"37a2", x"37a5", x"37a8", x"37ab", x"37ad", x"37b0", 
    x"37b3", x"37b6", x"37b9", x"37bc", x"37be", x"37c1", x"37c4", x"37c7", 
    x"37ca", x"37cd", x"37cf", x"37d2", x"37d5", x"37d8", x"37db", x"37de", 
    x"37e0", x"37e3", x"37e6", x"37e9", x"37ec", x"37ee", x"37f1", x"37f4", 
    x"37f7", x"37fa", x"37fd", x"37ff", x"3802", x"3805", x"3808", x"380b", 
    x"380e", x"3810", x"3813", x"3816", x"3819", x"381c", x"381e", x"3821", 
    x"3824", x"3827", x"382a", x"382d", x"382f", x"3832", x"3835", x"3838", 
    x"383b", x"383e", x"3840", x"3843", x"3846", x"3849", x"384c", x"384e", 
    x"3851", x"3854", x"3857", x"385a", x"385d", x"385f", x"3862", x"3865", 
    x"3868", x"386b", x"386d", x"3870", x"3873", x"3876", x"3879", x"387c", 
    x"387e", x"3881", x"3884", x"3887", x"388a", x"388d", x"388f", x"3892", 
    x"3895", x"3898", x"389b", x"389d", x"38a0", x"38a3", x"38a6", x"38a9", 
    x"38ab", x"38ae", x"38b1", x"38b4", x"38b7", x"38ba", x"38bc", x"38bf", 
    x"38c2", x"38c5", x"38c8", x"38ca", x"38cd", x"38d0", x"38d3", x"38d6", 
    x"38d9", x"38db", x"38de", x"38e1", x"38e4", x"38e7", x"38e9", x"38ec", 
    x"38ef", x"38f2", x"38f5", x"38f8", x"38fa", x"38fd", x"3900", x"3903", 
    x"3906", x"3908", x"390b", x"390e", x"3911", x"3914", x"3916", x"3919", 
    x"391c", x"391f", x"3922", x"3924", x"3927", x"392a", x"392d", x"3930", 
    x"3933", x"3935", x"3938", x"393b", x"393e", x"3941", x"3943", x"3946", 
    x"3949", x"394c", x"394f", x"3951", x"3954", x"3957", x"395a", x"395d", 
    x"3960", x"3962", x"3965", x"3968", x"396b", x"396e", x"3970", x"3973", 
    x"3976", x"3979", x"397c", x"397e", x"3981", x"3984", x"3987", x"398a", 
    x"398c", x"398f", x"3992", x"3995", x"3998", x"399a", x"399d", x"39a0", 
    x"39a3", x"39a6", x"39a8", x"39ab", x"39ae", x"39b1", x"39b4", x"39b6", 
    x"39b9", x"39bc", x"39bf", x"39c2", x"39c5", x"39c7", x"39ca", x"39cd", 
    x"39d0", x"39d3", x"39d5", x"39d8", x"39db", x"39de", x"39e1", x"39e3", 
    x"39e6", x"39e9", x"39ec", x"39ef", x"39f1", x"39f4", x"39f7", x"39fa", 
    x"39fd", x"39ff", x"3a02", x"3a05", x"3a08", x"3a0b", x"3a0d", x"3a10", 
    x"3a13", x"3a16", x"3a19", x"3a1b", x"3a1e", x"3a21", x"3a24", x"3a27", 
    x"3a29", x"3a2c", x"3a2f", x"3a32", x"3a35", x"3a37", x"3a3a", x"3a3d", 
    x"3a40", x"3a43", x"3a45", x"3a48", x"3a4b", x"3a4e", x"3a51", x"3a53", 
    x"3a56", x"3a59", x"3a5c", x"3a5e", x"3a61", x"3a64", x"3a67", x"3a6a", 
    x"3a6c", x"3a6f", x"3a72", x"3a75", x"3a78", x"3a7a", x"3a7d", x"3a80", 
    x"3a83", x"3a86", x"3a88", x"3a8b", x"3a8e", x"3a91", x"3a94", x"3a96", 
    x"3a99", x"3a9c", x"3a9f", x"3aa2", x"3aa4", x"3aa7", x"3aaa", x"3aad", 
    x"3ab0", x"3ab2", x"3ab5", x"3ab8", x"3abb", x"3abd", x"3ac0", x"3ac3", 
    x"3ac6", x"3ac9", x"3acb", x"3ace", x"3ad1", x"3ad4", x"3ad7", x"3ad9", 
    x"3adc", x"3adf", x"3ae2", x"3ae5", x"3ae7", x"3aea", x"3aed", x"3af0", 
    x"3af2", x"3af5", x"3af8", x"3afb", x"3afe", x"3b00", x"3b03", x"3b06", 
    x"3b09", x"3b0c", x"3b0e", x"3b11", x"3b14", x"3b17", x"3b19", x"3b1c", 
    x"3b1f", x"3b22", x"3b25", x"3b27", x"3b2a", x"3b2d", x"3b30", x"3b33", 
    x"3b35", x"3b38", x"3b3b", x"3b3e", x"3b40", x"3b43", x"3b46", x"3b49", 
    x"3b4c", x"3b4e", x"3b51", x"3b54", x"3b57", x"3b5a", x"3b5c", x"3b5f", 
    x"3b62", x"3b65", x"3b67", x"3b6a", x"3b6d", x"3b70", x"3b73", x"3b75", 
    x"3b78", x"3b7b", x"3b7e", x"3b81", x"3b83", x"3b86", x"3b89", x"3b8c", 
    x"3b8e", x"3b91", x"3b94", x"3b97", x"3b9a", x"3b9c", x"3b9f", x"3ba2", 
    x"3ba5", x"3ba7", x"3baa", x"3bad", x"3bb0", x"3bb3", x"3bb5", x"3bb8", 
    x"3bbb", x"3bbe", x"3bc0", x"3bc3", x"3bc6", x"3bc9", x"3bcc", x"3bce", 
    x"3bd1", x"3bd4", x"3bd7", x"3bd9", x"3bdc", x"3bdf", x"3be2", x"3be5", 
    x"3be7", x"3bea", x"3bed", x"3bf0", x"3bf2", x"3bf5", x"3bf8", x"3bfb", 
    x"3bfe", x"3c00", x"3c03", x"3c06", x"3c09", x"3c0b", x"3c0e", x"3c11", 
    x"3c14", x"3c16", x"3c19", x"3c1c", x"3c1f", x"3c22", x"3c24", x"3c27", 
    x"3c2a", x"3c2d", x"3c2f", x"3c32", x"3c35", x"3c38", x"3c3b", x"3c3d", 
    x"3c40", x"3c43", x"3c46", x"3c48", x"3c4b", x"3c4e", x"3c51", x"3c53", 
    x"3c56", x"3c59", x"3c5c", x"3c5f", x"3c61", x"3c64", x"3c67", x"3c6a", 
    x"3c6c", x"3c6f", x"3c72", x"3c75", x"3c77", x"3c7a", x"3c7d", x"3c80", 
    x"3c83", x"3c85", x"3c88", x"3c8b", x"3c8e", x"3c90", x"3c93", x"3c96", 
    x"3c99", x"3c9b", x"3c9e", x"3ca1", x"3ca4", x"3ca7", x"3ca9", x"3cac", 
    x"3caf", x"3cb2", x"3cb4", x"3cb7", x"3cba", x"3cbd", x"3cbf", x"3cc2", 
    x"3cc5", x"3cc8", x"3cca", x"3ccd", x"3cd0", x"3cd3", x"3cd6", x"3cd8", 
    x"3cdb", x"3cde", x"3ce1", x"3ce3", x"3ce6", x"3ce9", x"3cec", x"3cee", 
    x"3cf1", x"3cf4", x"3cf7", x"3cf9", x"3cfc", x"3cff", x"3d02", x"3d05", 
    x"3d07", x"3d0a", x"3d0d", x"3d10", x"3d12", x"3d15", x"3d18", x"3d1b", 
    x"3d1d", x"3d20", x"3d23", x"3d26", x"3d28", x"3d2b", x"3d2e", x"3d31", 
    x"3d33", x"3d36", x"3d39", x"3d3c", x"3d3e", x"3d41", x"3d44", x"3d47", 
    x"3d4a", x"3d4c", x"3d4f", x"3d52", x"3d55", x"3d57", x"3d5a", x"3d5d", 
    x"3d60", x"3d62", x"3d65", x"3d68", x"3d6b", x"3d6d", x"3d70", x"3d73", 
    x"3d76", x"3d78", x"3d7b", x"3d7e", x"3d81", x"3d83", x"3d86", x"3d89", 
    x"3d8c", x"3d8e", x"3d91", x"3d94", x"3d97", x"3d99", x"3d9c", x"3d9f", 
    x"3da2", x"3da4", x"3da7", x"3daa", x"3dad", x"3daf", x"3db2", x"3db5", 
    x"3db8", x"3dba", x"3dbd", x"3dc0", x"3dc3", x"3dc5", x"3dc8", x"3dcb", 
    x"3dce", x"3dd0", x"3dd3", x"3dd6", x"3dd9", x"3ddb", x"3dde", x"3de1", 
    x"3de4", x"3de6", x"3de9", x"3dec", x"3def", x"3df1", x"3df4", x"3df7", 
    x"3dfa", x"3dfc", x"3dff", x"3e02", x"3e05", x"3e07", x"3e0a", x"3e0d", 
    x"3e10", x"3e12", x"3e15", x"3e18", x"3e1b", x"3e1d", x"3e20", x"3e23", 
    x"3e26", x"3e28", x"3e2b", x"3e2e", x"3e31", x"3e33", x"3e36", x"3e39", 
    x"3e3c", x"3e3e", x"3e41", x"3e44", x"3e47", x"3e49", x"3e4c", x"3e4f", 
    x"3e52", x"3e54", x"3e57", x"3e5a", x"3e5d", x"3e5f", x"3e62", x"3e65", 
    x"3e68", x"3e6a", x"3e6d", x"3e70", x"3e73", x"3e75", x"3e78", x"3e7b", 
    x"3e7d", x"3e80", x"3e83", x"3e86", x"3e88", x"3e8b", x"3e8e", x"3e91", 
    x"3e93", x"3e96", x"3e99", x"3e9c", x"3e9e", x"3ea1", x"3ea4", x"3ea7", 
    x"3ea9", x"3eac", x"3eaf", x"3eb2", x"3eb4", x"3eb7", x"3eba", x"3ebd", 
    x"3ebf", x"3ec2", x"3ec5", x"3ec7", x"3eca", x"3ecd", x"3ed0", x"3ed2", 
    x"3ed5", x"3ed8", x"3edb", x"3edd", x"3ee0", x"3ee3", x"3ee6", x"3ee8", 
    x"3eeb", x"3eee", x"3ef1", x"3ef3", x"3ef6", x"3ef9", x"3efb", x"3efe", 
    x"3f01", x"3f04", x"3f06", x"3f09", x"3f0c", x"3f0f", x"3f11", x"3f14", 
    x"3f17", x"3f1a", x"3f1c", x"3f1f", x"3f22", x"3f24", x"3f27", x"3f2a", 
    x"3f2d", x"3f2f", x"3f32", x"3f35", x"3f38", x"3f3a", x"3f3d", x"3f40", 
    x"3f43", x"3f45", x"3f48", x"3f4b", x"3f4d", x"3f50", x"3f53", x"3f56", 
    x"3f58", x"3f5b", x"3f5e", x"3f61", x"3f63", x"3f66", x"3f69", x"3f6b", 
    x"3f6e", x"3f71", x"3f74", x"3f76", x"3f79", x"3f7c", x"3f7f", x"3f81", 
    x"3f84", x"3f87", x"3f89", x"3f8c", x"3f8f", x"3f92", x"3f94", x"3f97", 
    x"3f9a", x"3f9d", x"3f9f", x"3fa2", x"3fa5", x"3fa7", x"3faa", x"3fad", 
    x"3fb0", x"3fb2", x"3fb5", x"3fb8", x"3fbb", x"3fbd", x"3fc0", x"3fc3", 
    x"3fc5", x"3fc8", x"3fcb", x"3fce", x"3fd0", x"3fd3", x"3fd6", x"3fd8", 
    x"3fdb", x"3fde", x"3fe1", x"3fe3", x"3fe6", x"3fe9", x"3fec", x"3fee", 
    x"3ff1", x"3ff4", x"3ff6", x"3ff9", x"3ffc", x"3fff", x"4001", x"4004", 
    x"4007", x"4009", x"400c", x"400f", x"4012", x"4014", x"4017", x"401a", 
    x"401d", x"401f", x"4022", x"4025", x"4027", x"402a", x"402d", x"4030", 
    x"4032", x"4035", x"4038", x"403a", x"403d", x"4040", x"4043", x"4045", 
    x"4048", x"404b", x"404d", x"4050", x"4053", x"4056", x"4058", x"405b", 
    x"405e", x"4060", x"4063", x"4066", x"4069", x"406b", x"406e", x"4071", 
    x"4073", x"4076", x"4079", x"407c", x"407e", x"4081", x"4084", x"4086", 
    x"4089", x"408c", x"408f", x"4091", x"4094", x"4097", x"4099", x"409c", 
    x"409f", x"40a2", x"40a4", x"40a7", x"40aa", x"40ac", x"40af", x"40b2", 
    x"40b5", x"40b7", x"40ba", x"40bd", x"40bf", x"40c2", x"40c5", x"40c8", 
    x"40ca", x"40cd", x"40d0", x"40d2", x"40d5", x"40d8", x"40da", x"40dd", 
    x"40e0", x"40e3", x"40e5", x"40e8", x"40eb", x"40ed", x"40f0", x"40f3", 
    x"40f6", x"40f8", x"40fb", x"40fe", x"4100", x"4103", x"4106", x"4108", 
    x"410b", x"410e", x"4111", x"4113", x"4116", x"4119", x"411b", x"411e", 
    x"4121", x"4124", x"4126", x"4129", x"412c", x"412e", x"4131", x"4134", 
    x"4136", x"4139", x"413c", x"413f", x"4141", x"4144", x"4147", x"4149", 
    x"414c", x"414f", x"4151", x"4154", x"4157", x"415a", x"415c", x"415f", 
    x"4162", x"4164", x"4167", x"416a", x"416d", x"416f", x"4172", x"4175", 
    x"4177", x"417a", x"417d", x"417f", x"4182", x"4185", x"4187", x"418a", 
    x"418d", x"4190", x"4192", x"4195", x"4198", x"419a", x"419d", x"41a0", 
    x"41a2", x"41a5", x"41a8", x"41ab", x"41ad", x"41b0", x"41b3", x"41b5", 
    x"41b8", x"41bb", x"41bd", x"41c0", x"41c3", x"41c6", x"41c8", x"41cb", 
    x"41ce", x"41d0", x"41d3", x"41d6", x"41d8", x"41db", x"41de", x"41e0", 
    x"41e3", x"41e6", x"41e9", x"41eb", x"41ee", x"41f1", x"41f3", x"41f6", 
    x"41f9", x"41fb", x"41fe", x"4201", x"4203", x"4206", x"4209", x"420c", 
    x"420e", x"4211", x"4214", x"4216", x"4219", x"421c", x"421e", x"4221", 
    x"4224", x"4226", x"4229", x"422c", x"422f", x"4231", x"4234", x"4237", 
    x"4239", x"423c", x"423f", x"4241", x"4244", x"4247", x"4249", x"424c", 
    x"424f", x"4251", x"4254", x"4257", x"425a", x"425c", x"425f", x"4262", 
    x"4264", x"4267", x"426a", x"426c", x"426f", x"4272", x"4274", x"4277", 
    x"427a", x"427c", x"427f", x"4282", x"4284", x"4287", x"428a", x"428d", 
    x"428f", x"4292", x"4295", x"4297", x"429a", x"429d", x"429f", x"42a2", 
    x"42a5", x"42a7", x"42aa", x"42ad", x"42af", x"42b2", x"42b5", x"42b7", 
    x"42ba", x"42bd", x"42bf", x"42c2", x"42c5", x"42c8", x"42ca", x"42cd", 
    x"42d0", x"42d2", x"42d5", x"42d8", x"42da", x"42dd", x"42e0", x"42e2", 
    x"42e5", x"42e8", x"42ea", x"42ed", x"42f0", x"42f2", x"42f5", x"42f8", 
    x"42fa", x"42fd", x"4300", x"4302", x"4305", x"4308", x"430a", x"430d", 
    x"4310", x"4313", x"4315", x"4318", x"431b", x"431d", x"4320", x"4323", 
    x"4325", x"4328", x"432b", x"432d", x"4330", x"4333", x"4335", x"4338", 
    x"433b", x"433d", x"4340", x"4343", x"4345", x"4348", x"434b", x"434d", 
    x"4350", x"4353", x"4355", x"4358", x"435b", x"435d", x"4360", x"4363", 
    x"4365", x"4368", x"436b", x"436d", x"4370", x"4373", x"4375", x"4378", 
    x"437b", x"437d", x"4380", x"4383", x"4385", x"4388", x"438b", x"438d", 
    x"4390", x"4393", x"4395", x"4398", x"439b", x"439d", x"43a0", x"43a3", 
    x"43a5", x"43a8", x"43ab", x"43ad", x"43b0", x"43b3", x"43b5", x"43b8", 
    x"43bb", x"43bd", x"43c0", x"43c3", x"43c5", x"43c8", x"43cb", x"43cd", 
    x"43d0", x"43d3", x"43d5", x"43d8", x"43db", x"43dd", x"43e0", x"43e3", 
    x"43e5", x"43e8", x"43eb", x"43ed", x"43f0", x"43f3", x"43f5", x"43f8", 
    x"43fb", x"43fd", x"4400", x"4403", x"4405", x"4408", x"440b", x"440d", 
    x"4410", x"4413", x"4415", x"4418", x"441b", x"441d", x"4420", x"4423", 
    x"4425", x"4428", x"442b", x"442d", x"4430", x"4433", x"4435", x"4438", 
    x"443b", x"443d", x"4440", x"4442", x"4445", x"4448", x"444a", x"444d", 
    x"4450", x"4452", x"4455", x"4458", x"445a", x"445d", x"4460", x"4462", 
    x"4465", x"4468", x"446a", x"446d", x"4470", x"4472", x"4475", x"4478", 
    x"447a", x"447d", x"4480", x"4482", x"4485", x"4488", x"448a", x"448d", 
    x"448f", x"4492", x"4495", x"4497", x"449a", x"449d", x"449f", x"44a2", 
    x"44a5", x"44a7", x"44aa", x"44ad", x"44af", x"44b2", x"44b5", x"44b7", 
    x"44ba", x"44bd", x"44bf", x"44c2", x"44c5", x"44c7", x"44ca", x"44cc", 
    x"44cf", x"44d2", x"44d4", x"44d7", x"44da", x"44dc", x"44df", x"44e2", 
    x"44e4", x"44e7", x"44ea", x"44ec", x"44ef", x"44f2", x"44f4", x"44f7", 
    x"44f9", x"44fc", x"44ff", x"4501", x"4504", x"4507", x"4509", x"450c", 
    x"450f", x"4511", x"4514", x"4517", x"4519", x"451c", x"451f", x"4521", 
    x"4524", x"4526", x"4529", x"452c", x"452e", x"4531", x"4534", x"4536", 
    x"4539", x"453c", x"453e", x"4541", x"4544", x"4546", x"4549", x"454b", 
    x"454e", x"4551", x"4553", x"4556", x"4559", x"455b", x"455e", x"4561", 
    x"4563", x"4566", x"4568", x"456b", x"456e", x"4570", x"4573", x"4576", 
    x"4578", x"457b", x"457e", x"4580", x"4583", x"4586", x"4588", x"458b", 
    x"458d", x"4590", x"4593", x"4595", x"4598", x"459b", x"459d", x"45a0", 
    x"45a3", x"45a5", x"45a8", x"45aa", x"45ad", x"45b0", x"45b2", x"45b5", 
    x"45b8", x"45ba", x"45bd", x"45bf", x"45c2", x"45c5", x"45c7", x"45ca", 
    x"45cd", x"45cf", x"45d2", x"45d5", x"45d7", x"45da", x"45dc", x"45df", 
    x"45e2", x"45e4", x"45e7", x"45ea", x"45ec", x"45ef", x"45f2", x"45f4", 
    x"45f7", x"45f9", x"45fc", x"45ff", x"4601", x"4604", x"4607", x"4609", 
    x"460c", x"460e", x"4611", x"4614", x"4616", x"4619", x"461c", x"461e", 
    x"4621", x"4623", x"4626", x"4629", x"462b", x"462e", x"4631", x"4633", 
    x"4636", x"4638", x"463b", x"463e", x"4640", x"4643", x"4646", x"4648", 
    x"464b", x"464d", x"4650", x"4653", x"4655", x"4658", x"465b", x"465d", 
    x"4660", x"4662", x"4665", x"4668", x"466a", x"466d", x"4670", x"4672", 
    x"4675", x"4677", x"467a", x"467d", x"467f", x"4682", x"4685", x"4687", 
    x"468a", x"468c", x"468f", x"4692", x"4694", x"4697", x"469a", x"469c", 
    x"469f", x"46a1", x"46a4", x"46a7", x"46a9", x"46ac", x"46af", x"46b1", 
    x"46b4", x"46b6", x"46b9", x"46bc", x"46be", x"46c1", x"46c3", x"46c6", 
    x"46c9", x"46cb", x"46ce", x"46d1", x"46d3", x"46d6", x"46d8", x"46db", 
    x"46de", x"46e0", x"46e3", x"46e5", x"46e8", x"46eb", x"46ed", x"46f0", 
    x"46f3", x"46f5", x"46f8", x"46fa", x"46fd", x"4700", x"4702", x"4705", 
    x"4707", x"470a", x"470d", x"470f", x"4712", x"4715", x"4717", x"471a", 
    x"471c", x"471f", x"4722", x"4724", x"4727", x"4729", x"472c", x"472f", 
    x"4731", x"4734", x"4736", x"4739", x"473c", x"473e", x"4741", x"4744", 
    x"4746", x"4749", x"474b", x"474e", x"4751", x"4753", x"4756", x"4758", 
    x"475b", x"475e", x"4760", x"4763", x"4765", x"4768", x"476b", x"476d", 
    x"4770", x"4772", x"4775", x"4778", x"477a", x"477d", x"4780", x"4782", 
    x"4785", x"4787", x"478a", x"478d", x"478f", x"4792", x"4794", x"4797", 
    x"479a", x"479c", x"479f", x"47a1", x"47a4", x"47a7", x"47a9", x"47ac", 
    x"47ae", x"47b1", x"47b4", x"47b6", x"47b9", x"47bb", x"47be", x"47c1", 
    x"47c3", x"47c6", x"47c8", x"47cb", x"47ce", x"47d0", x"47d3", x"47d5", 
    x"47d8", x"47db", x"47dd", x"47e0", x"47e2", x"47e5", x"47e8", x"47ea", 
    x"47ed", x"47ef", x"47f2", x"47f5", x"47f7", x"47fa", x"47fc", x"47ff", 
    x"4802", x"4804", x"4807", x"4809", x"480c", x"480f", x"4811", x"4814", 
    x"4816", x"4819", x"481c", x"481e", x"4821", x"4823", x"4826", x"4829", 
    x"482b", x"482e", x"4830", x"4833", x"4835", x"4838", x"483b", x"483d", 
    x"4840", x"4842", x"4845", x"4848", x"484a", x"484d", x"484f", x"4852", 
    x"4855", x"4857", x"485a", x"485c", x"485f", x"4862", x"4864", x"4867", 
    x"4869", x"486c", x"486f", x"4871", x"4874", x"4876", x"4879", x"487b", 
    x"487e", x"4881", x"4883", x"4886", x"4888", x"488b", x"488e", x"4890", 
    x"4893", x"4895", x"4898", x"489b", x"489d", x"48a0", x"48a2", x"48a5", 
    x"48a7", x"48aa", x"48ad", x"48af", x"48b2", x"48b4", x"48b7", x"48ba", 
    x"48bc", x"48bf", x"48c1", x"48c4", x"48c6", x"48c9", x"48cc", x"48ce", 
    x"48d1", x"48d3", x"48d6", x"48d9", x"48db", x"48de", x"48e0", x"48e3", 
    x"48e5", x"48e8", x"48eb", x"48ed", x"48f0", x"48f2", x"48f5", x"48f8", 
    x"48fa", x"48fd", x"48ff", x"4902", x"4904", x"4907", x"490a", x"490c", 
    x"490f", x"4911", x"4914", x"4917", x"4919", x"491c", x"491e", x"4921", 
    x"4923", x"4926", x"4929", x"492b", x"492e", x"4930", x"4933", x"4935", 
    x"4938", x"493b", x"493d", x"4940", x"4942", x"4945", x"4947", x"494a", 
    x"494d", x"494f", x"4952", x"4954", x"4957", x"495a", x"495c", x"495f", 
    x"4961", x"4964", x"4966", x"4969", x"496c", x"496e", x"4971", x"4973", 
    x"4976", x"4978", x"497b", x"497e", x"4980", x"4983", x"4985", x"4988", 
    x"498a", x"498d", x"4990", x"4992", x"4995", x"4997", x"499a", x"499c", 
    x"499f", x"49a2", x"49a4", x"49a7", x"49a9", x"49ac", x"49ae", x"49b1", 
    x"49b4", x"49b6", x"49b9", x"49bb", x"49be", x"49c0", x"49c3", x"49c5", 
    x"49c8", x"49cb", x"49cd", x"49d0", x"49d2", x"49d5", x"49d7", x"49da", 
    x"49dd", x"49df", x"49e2", x"49e4", x"49e7", x"49e9", x"49ec", x"49ef", 
    x"49f1", x"49f4", x"49f6", x"49f9", x"49fb", x"49fe", x"4a00", x"4a03", 
    x"4a06", x"4a08", x"4a0b", x"4a0d", x"4a10", x"4a12", x"4a15", x"4a18", 
    x"4a1a", x"4a1d", x"4a1f", x"4a22", x"4a24", x"4a27", x"4a29", x"4a2c", 
    x"4a2f", x"4a31", x"4a34", x"4a36", x"4a39", x"4a3b", x"4a3e", x"4a41", 
    x"4a43", x"4a46", x"4a48", x"4a4b", x"4a4d", x"4a50", x"4a52", x"4a55", 
    x"4a58", x"4a5a", x"4a5d", x"4a5f", x"4a62", x"4a64", x"4a67", x"4a69", 
    x"4a6c", x"4a6f", x"4a71", x"4a74", x"4a76", x"4a79", x"4a7b", x"4a7e", 
    x"4a80", x"4a83", x"4a86", x"4a88", x"4a8b", x"4a8d", x"4a90", x"4a92", 
    x"4a95", x"4a97", x"4a9a", x"4a9d", x"4a9f", x"4aa2", x"4aa4", x"4aa7", 
    x"4aa9", x"4aac", x"4aae", x"4ab1", x"4ab3", x"4ab6", x"4ab9", x"4abb", 
    x"4abe", x"4ac0", x"4ac3", x"4ac5", x"4ac8", x"4aca", x"4acd", x"4ad0", 
    x"4ad2", x"4ad5", x"4ad7", x"4ada", x"4adc", x"4adf", x"4ae1", x"4ae4", 
    x"4ae6", x"4ae9", x"4aec", x"4aee", x"4af1", x"4af3", x"4af6", x"4af8", 
    x"4afb", x"4afd", x"4b00", x"4b02", x"4b05", x"4b08", x"4b0a", x"4b0d", 
    x"4b0f", x"4b12", x"4b14", x"4b17", x"4b19", x"4b1c", x"4b1e", x"4b21", 
    x"4b24", x"4b26", x"4b29", x"4b2b", x"4b2e", x"4b30", x"4b33", x"4b35", 
    x"4b38", x"4b3a", x"4b3d", x"4b40", x"4b42", x"4b45", x"4b47", x"4b4a", 
    x"4b4c", x"4b4f", x"4b51", x"4b54", x"4b56", x"4b59", x"4b5b", x"4b5e", 
    x"4b61", x"4b63", x"4b66", x"4b68", x"4b6b", x"4b6d", x"4b70", x"4b72", 
    x"4b75", x"4b77", x"4b7a", x"4b7c", x"4b7f", x"4b82", x"4b84", x"4b87", 
    x"4b89", x"4b8c", x"4b8e", x"4b91", x"4b93", x"4b96", x"4b98", x"4b9b", 
    x"4b9d", x"4ba0", x"4ba2", x"4ba5", x"4ba8", x"4baa", x"4bad", x"4baf", 
    x"4bb2", x"4bb4", x"4bb7", x"4bb9", x"4bbc", x"4bbe", x"4bc1", x"4bc3", 
    x"4bc6", x"4bc8", x"4bcb", x"4bce", x"4bd0", x"4bd3", x"4bd5", x"4bd8", 
    x"4bda", x"4bdd", x"4bdf", x"4be2", x"4be4", x"4be7", x"4be9", x"4bec", 
    x"4bee", x"4bf1", x"4bf4", x"4bf6", x"4bf9", x"4bfb", x"4bfe", x"4c00", 
    x"4c03", x"4c05", x"4c08", x"4c0a", x"4c0d", x"4c0f", x"4c12", x"4c14", 
    x"4c17", x"4c19", x"4c1c", x"4c1e", x"4c21", x"4c24", x"4c26", x"4c29", 
    x"4c2b", x"4c2e", x"4c30", x"4c33", x"4c35", x"4c38", x"4c3a", x"4c3d", 
    x"4c3f", x"4c42", x"4c44", x"4c47", x"4c49", x"4c4c", x"4c4e", x"4c51", 
    x"4c53", x"4c56", x"4c59", x"4c5b", x"4c5e", x"4c60", x"4c63", x"4c65", 
    x"4c68", x"4c6a", x"4c6d", x"4c6f", x"4c72", x"4c74", x"4c77", x"4c79", 
    x"4c7c", x"4c7e", x"4c81", x"4c83", x"4c86", x"4c88", x"4c8b", x"4c8d", 
    x"4c90", x"4c92", x"4c95", x"4c97", x"4c9a", x"4c9d", x"4c9f", x"4ca2", 
    x"4ca4", x"4ca7", x"4ca9", x"4cac", x"4cae", x"4cb1", x"4cb3", x"4cb6", 
    x"4cb8", x"4cbb", x"4cbd", x"4cc0", x"4cc2", x"4cc5", x"4cc7", x"4cca", 
    x"4ccc", x"4ccf", x"4cd1", x"4cd4", x"4cd6", x"4cd9", x"4cdb", x"4cde", 
    x"4ce0", x"4ce3", x"4ce5", x"4ce8", x"4cea", x"4ced", x"4cef", x"4cf2", 
    x"4cf4", x"4cf7", x"4cfa", x"4cfc", x"4cff", x"4d01", x"4d04", x"4d06", 
    x"4d09", x"4d0b", x"4d0e", x"4d10", x"4d13", x"4d15", x"4d18", x"4d1a", 
    x"4d1d", x"4d1f", x"4d22", x"4d24", x"4d27", x"4d29", x"4d2c", x"4d2e", 
    x"4d31", x"4d33", x"4d36", x"4d38", x"4d3b", x"4d3d", x"4d40", x"4d42", 
    x"4d45", x"4d47", x"4d4a", x"4d4c", x"4d4f", x"4d51", x"4d54", x"4d56", 
    x"4d59", x"4d5b", x"4d5e", x"4d60", x"4d63", x"4d65", x"4d68", x"4d6a", 
    x"4d6d", x"4d6f", x"4d72", x"4d74", x"4d77", x"4d79", x"4d7c", x"4d7e", 
    x"4d81", x"4d83", x"4d86", x"4d88", x"4d8b", x"4d8d", x"4d90", x"4d92", 
    x"4d95", x"4d97", x"4d9a", x"4d9c", x"4d9f", x"4da1", x"4da4", x"4da6", 
    x"4da9", x"4dab", x"4dae", x"4db0", x"4db3", x"4db5", x"4db8", x"4dba", 
    x"4dbd", x"4dbf", x"4dc2", x"4dc4", x"4dc7", x"4dc9", x"4dcc", x"4dce", 
    x"4dd1", x"4dd3", x"4dd6", x"4dd8", x"4ddb", x"4ddd", x"4de0", x"4de2", 
    x"4de5", x"4de7", x"4dea", x"4dec", x"4def", x"4df1", x"4df4", x"4df6", 
    x"4df9", x"4dfb", x"4dfe", x"4e00", x"4e03", x"4e05", x"4e08", x"4e0a", 
    x"4e0d", x"4e0f", x"4e11", x"4e14", x"4e16", x"4e19", x"4e1b", x"4e1e", 
    x"4e20", x"4e23", x"4e25", x"4e28", x"4e2a", x"4e2d", x"4e2f", x"4e32", 
    x"4e34", x"4e37", x"4e39", x"4e3c", x"4e3e", x"4e41", x"4e43", x"4e46", 
    x"4e48", x"4e4b", x"4e4d", x"4e50", x"4e52", x"4e55", x"4e57", x"4e5a", 
    x"4e5c", x"4e5f", x"4e61", x"4e64", x"4e66", x"4e68", x"4e6b", x"4e6d", 
    x"4e70", x"4e72", x"4e75", x"4e77", x"4e7a", x"4e7c", x"4e7f", x"4e81", 
    x"4e84", x"4e86", x"4e89", x"4e8b", x"4e8e", x"4e90", x"4e93", x"4e95", 
    x"4e98", x"4e9a", x"4e9d", x"4e9f", x"4ea2", x"4ea4", x"4ea7", x"4ea9", 
    x"4eab", x"4eae", x"4eb0", x"4eb3", x"4eb5", x"4eb8", x"4eba", x"4ebd", 
    x"4ebf", x"4ec2", x"4ec4", x"4ec7", x"4ec9", x"4ecc", x"4ece", x"4ed1", 
    x"4ed3", x"4ed6", x"4ed8", x"4edb", x"4edd", x"4edf", x"4ee2", x"4ee4", 
    x"4ee7", x"4ee9", x"4eec", x"4eee", x"4ef1", x"4ef3", x"4ef6", x"4ef8", 
    x"4efb", x"4efd", x"4f00", x"4f02", x"4f05", x"4f07", x"4f0a", x"4f0c", 
    x"4f0e", x"4f11", x"4f13", x"4f16", x"4f18", x"4f1b", x"4f1d", x"4f20", 
    x"4f22", x"4f25", x"4f27", x"4f2a", x"4f2c", x"4f2f", x"4f31", x"4f33", 
    x"4f36", x"4f38", x"4f3b", x"4f3d", x"4f40", x"4f42", x"4f45", x"4f47", 
    x"4f4a", x"4f4c", x"4f4f", x"4f51", x"4f54", x"4f56", x"4f58", x"4f5b", 
    x"4f5d", x"4f60", x"4f62", x"4f65", x"4f67", x"4f6a", x"4f6c", x"4f6f", 
    x"4f71", x"4f74", x"4f76", x"4f79", x"4f7b", x"4f7d", x"4f80", x"4f82", 
    x"4f85", x"4f87", x"4f8a", x"4f8c", x"4f8f", x"4f91", x"4f94", x"4f96", 
    x"4f99", x"4f9b", x"4f9d", x"4fa0", x"4fa2", x"4fa5", x"4fa7", x"4faa", 
    x"4fac", x"4faf", x"4fb1", x"4fb4", x"4fb6", x"4fb8", x"4fbb", x"4fbd", 
    x"4fc0", x"4fc2", x"4fc5", x"4fc7", x"4fca", x"4fcc", x"4fcf", x"4fd1", 
    x"4fd4", x"4fd6", x"4fd8", x"4fdb", x"4fdd", x"4fe0", x"4fe2", x"4fe5", 
    x"4fe7", x"4fea", x"4fec", x"4fef", x"4ff1", x"4ff3", x"4ff6", x"4ff8", 
    x"4ffb", x"4ffd", x"5000", x"5002", x"5005", x"5007", x"5009", x"500c", 
    x"500e", x"5011", x"5013", x"5016", x"5018", x"501b", x"501d", x"5020", 
    x"5022", x"5024", x"5027", x"5029", x"502c", x"502e", x"5031", x"5033", 
    x"5036", x"5038", x"503a", x"503d", x"503f", x"5042", x"5044", x"5047", 
    x"5049", x"504c", x"504e", x"5050", x"5053", x"5055", x"5058", x"505a", 
    x"505d", x"505f", x"5062", x"5064", x"5067", x"5069", x"506b", x"506e", 
    x"5070", x"5073", x"5075", x"5078", x"507a", x"507c", x"507f", x"5081", 
    x"5084", x"5086", x"5089", x"508b", x"508e", x"5090", x"5092", x"5095", 
    x"5097", x"509a", x"509c", x"509f", x"50a1", x"50a4", x"50a6", x"50a8", 
    x"50ab", x"50ad", x"50b0", x"50b2", x"50b5", x"50b7", x"50ba", x"50bc", 
    x"50be", x"50c1", x"50c3", x"50c6", x"50c8", x"50cb", x"50cd", x"50cf", 
    x"50d2", x"50d4", x"50d7", x"50d9", x"50dc", x"50de", x"50e0", x"50e3", 
    x"50e5", x"50e8", x"50ea", x"50ed", x"50ef", x"50f2", x"50f4", x"50f6", 
    x"50f9", x"50fb", x"50fe", x"5100", x"5103", x"5105", x"5107", x"510a", 
    x"510c", x"510f", x"5111", x"5114", x"5116", x"5118", x"511b", x"511d", 
    x"5120", x"5122", x"5125", x"5127", x"5129", x"512c", x"512e", x"5131", 
    x"5133", x"5136", x"5138", x"513a", x"513d", x"513f", x"5142", x"5144", 
    x"5147", x"5149", x"514b", x"514e", x"5150", x"5153", x"5155", x"5158", 
    x"515a", x"515c", x"515f", x"5161", x"5164", x"5166", x"5169", x"516b", 
    x"516d", x"5170", x"5172", x"5175", x"5177", x"517a", x"517c", x"517e", 
    x"5181", x"5183", x"5186", x"5188", x"518a", x"518d", x"518f", x"5192", 
    x"5194", x"5197", x"5199", x"519b", x"519e", x"51a0", x"51a3", x"51a5", 
    x"51a8", x"51aa", x"51ac", x"51af", x"51b1", x"51b4", x"51b6", x"51b8", 
    x"51bb", x"51bd", x"51c0", x"51c2", x"51c5", x"51c7", x"51c9", x"51cc", 
    x"51ce", x"51d1", x"51d3", x"51d5", x"51d8", x"51da", x"51dd", x"51df", 
    x"51e2", x"51e4", x"51e6", x"51e9", x"51eb", x"51ee", x"51f0", x"51f2", 
    x"51f5", x"51f7", x"51fa", x"51fc", x"51fe", x"5201", x"5203", x"5206", 
    x"5208", x"520b", x"520d", x"520f", x"5212", x"5214", x"5217", x"5219", 
    x"521b", x"521e", x"5220", x"5223", x"5225", x"5227", x"522a", x"522c", 
    x"522f", x"5231", x"5233", x"5236", x"5238", x"523b", x"523d", x"5240", 
    x"5242", x"5244", x"5247", x"5249", x"524c", x"524e", x"5250", x"5253", 
    x"5255", x"5258", x"525a", x"525c", x"525f", x"5261", x"5264", x"5266", 
    x"5268", x"526b", x"526d", x"5270", x"5272", x"5274", x"5277", x"5279", 
    x"527c", x"527e", x"5280", x"5283", x"5285", x"5288", x"528a", x"528c", 
    x"528f", x"5291", x"5294", x"5296", x"5298", x"529b", x"529d", x"52a0", 
    x"52a2", x"52a4", x"52a7", x"52a9", x"52ac", x"52ae", x"52b0", x"52b3", 
    x"52b5", x"52b8", x"52ba", x"52bc", x"52bf", x"52c1", x"52c4", x"52c6", 
    x"52c8", x"52cb", x"52cd", x"52d0", x"52d2", x"52d4", x"52d7", x"52d9", 
    x"52dc", x"52de", x"52e0", x"52e3", x"52e5", x"52e8", x"52ea", x"52ec", 
    x"52ef", x"52f1", x"52f4", x"52f6", x"52f8", x"52fb", x"52fd", x"52ff", 
    x"5302", x"5304", x"5307", x"5309", x"530b", x"530e", x"5310", x"5313", 
    x"5315", x"5317", x"531a", x"531c", x"531f", x"5321", x"5323", x"5326", 
    x"5328", x"532a", x"532d", x"532f", x"5332", x"5334", x"5336", x"5339", 
    x"533b", x"533e", x"5340", x"5342", x"5345", x"5347", x"534a", x"534c", 
    x"534e", x"5351", x"5353", x"5355", x"5358", x"535a", x"535d", x"535f", 
    x"5361", x"5364", x"5366", x"5369", x"536b", x"536d", x"5370", x"5372", 
    x"5374", x"5377", x"5379", x"537c", x"537e", x"5380", x"5383", x"5385", 
    x"5387", x"538a", x"538c", x"538f", x"5391", x"5393", x"5396", x"5398", 
    x"539b", x"539d", x"539f", x"53a2", x"53a4", x"53a6", x"53a9", x"53ab", 
    x"53ae", x"53b0", x"53b2", x"53b5", x"53b7", x"53b9", x"53bc", x"53be", 
    x"53c1", x"53c3", x"53c5", x"53c8", x"53ca", x"53cc", x"53cf", x"53d1", 
    x"53d4", x"53d6", x"53d8", x"53db", x"53dd", x"53df", x"53e2", x"53e4", 
    x"53e7", x"53e9", x"53eb", x"53ee", x"53f0", x"53f2", x"53f5", x"53f7", 
    x"53fa", x"53fc", x"53fe", x"5401", x"5403", x"5405", x"5408", x"540a", 
    x"540c", x"540f", x"5411", x"5414", x"5416", x"5418", x"541b", x"541d", 
    x"541f", x"5422", x"5424", x"5427", x"5429", x"542b", x"542e", x"5430", 
    x"5432", x"5435", x"5437", x"5439", x"543c", x"543e", x"5441", x"5443", 
    x"5445", x"5448", x"544a", x"544c", x"544f", x"5451", x"5453", x"5456", 
    x"5458", x"545b", x"545d", x"545f", x"5462", x"5464", x"5466", x"5469", 
    x"546b", x"546d", x"5470", x"5472", x"5475", x"5477", x"5479", x"547c", 
    x"547e", x"5480", x"5483", x"5485", x"5487", x"548a", x"548c", x"548e", 
    x"5491", x"5493", x"5496", x"5498", x"549a", x"549d", x"549f", x"54a1", 
    x"54a4", x"54a6", x"54a8", x"54ab", x"54ad", x"54af", x"54b2", x"54b4", 
    x"54b7", x"54b9", x"54bb", x"54be", x"54c0", x"54c2", x"54c5", x"54c7", 
    x"54c9", x"54cc", x"54ce", x"54d0", x"54d3", x"54d5", x"54d7", x"54da", 
    x"54dc", x"54df", x"54e1", x"54e3", x"54e6", x"54e8", x"54ea", x"54ed", 
    x"54ef", x"54f1", x"54f4", x"54f6", x"54f8", x"54fb", x"54fd", x"54ff", 
    x"5502", x"5504", x"5506", x"5509", x"550b", x"550e", x"5510", x"5512", 
    x"5515", x"5517", x"5519", x"551c", x"551e", x"5520", x"5523", x"5525", 
    x"5527", x"552a", x"552c", x"552e", x"5531", x"5533", x"5535", x"5538", 
    x"553a", x"553c", x"553f", x"5541", x"5543", x"5546", x"5548", x"554b", 
    x"554d", x"554f", x"5552", x"5554", x"5556", x"5559", x"555b", x"555d", 
    x"5560", x"5562", x"5564", x"5567", x"5569", x"556b", x"556e", x"5570", 
    x"5572", x"5575", x"5577", x"5579", x"557c", x"557e", x"5580", x"5583", 
    x"5585", x"5587", x"558a", x"558c", x"558e", x"5591", x"5593", x"5595", 
    x"5598", x"559a", x"559c", x"559f", x"55a1", x"55a3", x"55a6", x"55a8", 
    x"55aa", x"55ad", x"55af", x"55b1", x"55b4", x"55b6", x"55b8", x"55bb", 
    x"55bd", x"55bf", x"55c2", x"55c4", x"55c6", x"55c9", x"55cb", x"55cd", 
    x"55d0", x"55d2", x"55d4", x"55d7", x"55d9", x"55db", x"55de", x"55e0", 
    x"55e2", x"55e5", x"55e7", x"55e9", x"55ec", x"55ee", x"55f0", x"55f3", 
    x"55f5", x"55f7", x"55fa", x"55fc", x"55fe", x"5601", x"5603", x"5605", 
    x"5608", x"560a", x"560c", x"560f", x"5611", x"5613", x"5616", x"5618", 
    x"561a", x"561d", x"561f", x"5621", x"5623", x"5626", x"5628", x"562a", 
    x"562d", x"562f", x"5631", x"5634", x"5636", x"5638", x"563b", x"563d", 
    x"563f", x"5642", x"5644", x"5646", x"5649", x"564b", x"564d", x"5650", 
    x"5652", x"5654", x"5657", x"5659", x"565b", x"565e", x"5660", x"5662", 
    x"5664", x"5667", x"5669", x"566b", x"566e", x"5670", x"5672", x"5675", 
    x"5677", x"5679", x"567c", x"567e", x"5680", x"5683", x"5685", x"5687", 
    x"568a", x"568c", x"568e", x"5690", x"5693", x"5695", x"5697", x"569a", 
    x"569c", x"569e", x"56a1", x"56a3", x"56a5", x"56a8", x"56aa", x"56ac", 
    x"56af", x"56b1", x"56b3", x"56b5", x"56b8", x"56ba", x"56bc", x"56bf", 
    x"56c1", x"56c3", x"56c6", x"56c8", x"56ca", x"56cd", x"56cf", x"56d1", 
    x"56d3", x"56d6", x"56d8", x"56da", x"56dd", x"56df", x"56e1", x"56e4", 
    x"56e6", x"56e8", x"56eb", x"56ed", x"56ef", x"56f1", x"56f4", x"56f6", 
    x"56f8", x"56fb", x"56fd", x"56ff", x"5702", x"5704", x"5706", x"5709", 
    x"570b", x"570d", x"570f", x"5712", x"5714", x"5716", x"5719", x"571b", 
    x"571d", x"5720", x"5722", x"5724", x"5726", x"5729", x"572b", x"572d", 
    x"5730", x"5732", x"5734", x"5737", x"5739", x"573b", x"573d", x"5740", 
    x"5742", x"5744", x"5747", x"5749", x"574b", x"574e", x"5750", x"5752", 
    x"5754", x"5757", x"5759", x"575b", x"575e", x"5760", x"5762", x"5765", 
    x"5767", x"5769", x"576b", x"576e", x"5770", x"5772", x"5775", x"5777", 
    x"5779", x"577b", x"577e", x"5780", x"5782", x"5785", x"5787", x"5789", 
    x"578b", x"578e", x"5790", x"5792", x"5795", x"5797", x"5799", x"579c", 
    x"579e", x"57a0", x"57a2", x"57a5", x"57a7", x"57a9", x"57ac", x"57ae", 
    x"57b0", x"57b2", x"57b5", x"57b7", x"57b9", x"57bc", x"57be", x"57c0", 
    x"57c2", x"57c5", x"57c7", x"57c9", x"57cc", x"57ce", x"57d0", x"57d2", 
    x"57d5", x"57d7", x"57d9", x"57dc", x"57de", x"57e0", x"57e2", x"57e5", 
    x"57e7", x"57e9", x"57ec", x"57ee", x"57f0", x"57f2", x"57f5", x"57f7", 
    x"57f9", x"57fc", x"57fe", x"5800", x"5802", x"5805", x"5807", x"5809", 
    x"580c", x"580e", x"5810", x"5812", x"5815", x"5817", x"5819", x"581b", 
    x"581e", x"5820", x"5822", x"5825", x"5827", x"5829", x"582b", x"582e", 
    x"5830", x"5832", x"5835", x"5837", x"5839", x"583b", x"583e", x"5840", 
    x"5842", x"5844", x"5847", x"5849", x"584b", x"584e", x"5850", x"5852", 
    x"5854", x"5857", x"5859", x"585b", x"585d", x"5860", x"5862", x"5864", 
    x"5867", x"5869", x"586b", x"586d", x"5870", x"5872", x"5874", x"5876", 
    x"5879", x"587b", x"587d", x"5880", x"5882", x"5884", x"5886", x"5889", 
    x"588b", x"588d", x"588f", x"5892", x"5894", x"5896", x"5898", x"589b", 
    x"589d", x"589f", x"58a2", x"58a4", x"58a6", x"58a8", x"58ab", x"58ad", 
    x"58af", x"58b1", x"58b4", x"58b6", x"58b8", x"58ba", x"58bd", x"58bf", 
    x"58c1", x"58c4", x"58c6", x"58c8", x"58ca", x"58cd", x"58cf", x"58d1", 
    x"58d3", x"58d6", x"58d8", x"58da", x"58dc", x"58df", x"58e1", x"58e3", 
    x"58e5", x"58e8", x"58ea", x"58ec", x"58ee", x"58f1", x"58f3", x"58f5", 
    x"58f8", x"58fa", x"58fc", x"58fe", x"5901", x"5903", x"5905", x"5907", 
    x"590a", x"590c", x"590e", x"5910", x"5913", x"5915", x"5917", x"5919", 
    x"591c", x"591e", x"5920", x"5922", x"5925", x"5927", x"5929", x"592b", 
    x"592e", x"5930", x"5932", x"5934", x"5937", x"5939", x"593b", x"593d", 
    x"5940", x"5942", x"5944", x"5946", x"5949", x"594b", x"594d", x"594f", 
    x"5952", x"5954", x"5956", x"5958", x"595b", x"595d", x"595f", x"5961", 
    x"5964", x"5966", x"5968", x"596a", x"596d", x"596f", x"5971", x"5973", 
    x"5976", x"5978", x"597a", x"597c", x"597f", x"5981", x"5983", x"5985", 
    x"5988", x"598a", x"598c", x"598e", x"5991", x"5993", x"5995", x"5997", 
    x"599a", x"599c", x"599e", x"59a0", x"59a3", x"59a5", x"59a7", x"59a9", 
    x"59ac", x"59ae", x"59b0", x"59b2", x"59b5", x"59b7", x"59b9", x"59bb", 
    x"59bd", x"59c0", x"59c2", x"59c4", x"59c6", x"59c9", x"59cb", x"59cd", 
    x"59cf", x"59d2", x"59d4", x"59d6", x"59d8", x"59db", x"59dd", x"59df", 
    x"59e1", x"59e4", x"59e6", x"59e8", x"59ea", x"59ec", x"59ef", x"59f1", 
    x"59f3", x"59f5", x"59f8", x"59fa", x"59fc", x"59fe", x"5a01", x"5a03", 
    x"5a05", x"5a07", x"5a0a", x"5a0c", x"5a0e", x"5a10", x"5a12", x"5a15", 
    x"5a17", x"5a19", x"5a1b", x"5a1e", x"5a20", x"5a22", x"5a24", x"5a27", 
    x"5a29", x"5a2b", x"5a2d", x"5a2f", x"5a32", x"5a34", x"5a36", x"5a38", 
    x"5a3b", x"5a3d", x"5a3f", x"5a41", x"5a43", x"5a46", x"5a48", x"5a4a", 
    x"5a4c", x"5a4f", x"5a51", x"5a53", x"5a55", x"5a58", x"5a5a", x"5a5c", 
    x"5a5e", x"5a60", x"5a63", x"5a65", x"5a67", x"5a69", x"5a6c", x"5a6e", 
    x"5a70", x"5a72", x"5a74", x"5a77", x"5a79", x"5a7b", x"5a7d", x"5a80", 
    x"5a82", x"5a84", x"5a86", x"5a88", x"5a8b", x"5a8d", x"5a8f", x"5a91", 
    x"5a94", x"5a96", x"5a98", x"5a9a", x"5a9c", x"5a9f", x"5aa1", x"5aa3", 
    x"5aa5", x"5aa8", x"5aaa", x"5aac", x"5aae", x"5ab0", x"5ab3", x"5ab5", 
    x"5ab7", x"5ab9", x"5abb", x"5abe", x"5ac0", x"5ac2", x"5ac4", x"5ac7", 
    x"5ac9", x"5acb", x"5acd", x"5acf", x"5ad2", x"5ad4", x"5ad6", x"5ad8", 
    x"5ada", x"5add", x"5adf", x"5ae1", x"5ae3", x"5ae6", x"5ae8", x"5aea", 
    x"5aec", x"5aee", x"5af1", x"5af3", x"5af5", x"5af7", x"5af9", x"5afc", 
    x"5afe", x"5b00", x"5b02", x"5b04", x"5b07", x"5b09", x"5b0b", x"5b0d", 
    x"5b0f", x"5b12", x"5b14", x"5b16", x"5b18", x"5b1b", x"5b1d", x"5b1f", 
    x"5b21", x"5b23", x"5b26", x"5b28", x"5b2a", x"5b2c", x"5b2e", x"5b31", 
    x"5b33", x"5b35", x"5b37", x"5b39", x"5b3c", x"5b3e", x"5b40", x"5b42", 
    x"5b44", x"5b47", x"5b49", x"5b4b", x"5b4d", x"5b4f", x"5b52", x"5b54", 
    x"5b56", x"5b58", x"5b5a", x"5b5d", x"5b5f", x"5b61", x"5b63", x"5b65", 
    x"5b68", x"5b6a", x"5b6c", x"5b6e", x"5b70", x"5b73", x"5b75", x"5b77", 
    x"5b79", x"5b7b", x"5b7e", x"5b80", x"5b82", x"5b84", x"5b86", x"5b89", 
    x"5b8b", x"5b8d", x"5b8f", x"5b91", x"5b94", x"5b96", x"5b98", x"5b9a", 
    x"5b9c", x"5b9f", x"5ba1", x"5ba3", x"5ba5", x"5ba7", x"5baa", x"5bac", 
    x"5bae", x"5bb0", x"5bb2", x"5bb4", x"5bb7", x"5bb9", x"5bbb", x"5bbd", 
    x"5bbf", x"5bc2", x"5bc4", x"5bc6", x"5bc8", x"5bca", x"5bcd", x"5bcf", 
    x"5bd1", x"5bd3", x"5bd5", x"5bd8", x"5bda", x"5bdc", x"5bde", x"5be0", 
    x"5be2", x"5be5", x"5be7", x"5be9", x"5beb", x"5bed", x"5bf0", x"5bf2", 
    x"5bf4", x"5bf6", x"5bf8", x"5bfa", x"5bfd", x"5bff", x"5c01", x"5c03", 
    x"5c05", x"5c08", x"5c0a", x"5c0c", x"5c0e", x"5c10", x"5c13", x"5c15", 
    x"5c17", x"5c19", x"5c1b", x"5c1d", x"5c20", x"5c22", x"5c24", x"5c26", 
    x"5c28", x"5c2b", x"5c2d", x"5c2f", x"5c31", x"5c33", x"5c35", x"5c38", 
    x"5c3a", x"5c3c", x"5c3e", x"5c40", x"5c42", x"5c45", x"5c47", x"5c49", 
    x"5c4b", x"5c4d", x"5c50", x"5c52", x"5c54", x"5c56", x"5c58", x"5c5a", 
    x"5c5d", x"5c5f", x"5c61", x"5c63", x"5c65", x"5c67", x"5c6a", x"5c6c", 
    x"5c6e", x"5c70", x"5c72", x"5c74", x"5c77", x"5c79", x"5c7b", x"5c7d", 
    x"5c7f", x"5c82", x"5c84", x"5c86", x"5c88", x"5c8a", x"5c8c", x"5c8f", 
    x"5c91", x"5c93", x"5c95", x"5c97", x"5c99", x"5c9c", x"5c9e", x"5ca0", 
    x"5ca2", x"5ca4", x"5ca6", x"5ca9", x"5cab", x"5cad", x"5caf", x"5cb1", 
    x"5cb3", x"5cb6", x"5cb8", x"5cba", x"5cbc", x"5cbe", x"5cc0", x"5cc3", 
    x"5cc5", x"5cc7", x"5cc9", x"5ccb", x"5ccd", x"5cd0", x"5cd2", x"5cd4", 
    x"5cd6", x"5cd8", x"5cda", x"5cdd", x"5cdf", x"5ce1", x"5ce3", x"5ce5", 
    x"5ce7", x"5ce9", x"5cec", x"5cee", x"5cf0", x"5cf2", x"5cf4", x"5cf6", 
    x"5cf9", x"5cfb", x"5cfd", x"5cff", x"5d01", x"5d03", x"5d06", x"5d08", 
    x"5d0a", x"5d0c", x"5d0e", x"5d10", x"5d13", x"5d15", x"5d17", x"5d19", 
    x"5d1b", x"5d1d", x"5d1f", x"5d22", x"5d24", x"5d26", x"5d28", x"5d2a", 
    x"5d2c", x"5d2f", x"5d31", x"5d33", x"5d35", x"5d37", x"5d39", x"5d3b", 
    x"5d3e", x"5d40", x"5d42", x"5d44", x"5d46", x"5d48", x"5d4b", x"5d4d", 
    x"5d4f", x"5d51", x"5d53", x"5d55", x"5d57", x"5d5a", x"5d5c", x"5d5e", 
    x"5d60", x"5d62", x"5d64", x"5d66", x"5d69", x"5d6b", x"5d6d", x"5d6f", 
    x"5d71", x"5d73", x"5d75", x"5d78", x"5d7a", x"5d7c", x"5d7e", x"5d80", 
    x"5d82", x"5d84", x"5d87", x"5d89", x"5d8b", x"5d8d", x"5d8f", x"5d91", 
    x"5d94", x"5d96", x"5d98", x"5d9a", x"5d9c", x"5d9e", x"5da0", x"5da3", 
    x"5da5", x"5da7", x"5da9", x"5dab", x"5dad", x"5daf", x"5db1", x"5db4", 
    x"5db6", x"5db8", x"5dba", x"5dbc", x"5dbe", x"5dc0", x"5dc3", x"5dc5", 
    x"5dc7", x"5dc9", x"5dcb", x"5dcd", x"5dcf", x"5dd2", x"5dd4", x"5dd6", 
    x"5dd8", x"5dda", x"5ddc", x"5dde", x"5de1", x"5de3", x"5de5", x"5de7", 
    x"5de9", x"5deb", x"5ded", x"5def", x"5df2", x"5df4", x"5df6", x"5df8", 
    x"5dfa", x"5dfc", x"5dfe", x"5e01", x"5e03", x"5e05", x"5e07", x"5e09", 
    x"5e0b", x"5e0d", x"5e0f", x"5e12", x"5e14", x"5e16", x"5e18", x"5e1a", 
    x"5e1c", x"5e1e", x"5e20", x"5e23", x"5e25", x"5e27", x"5e29", x"5e2b", 
    x"5e2d", x"5e2f", x"5e32", x"5e34", x"5e36", x"5e38", x"5e3a", x"5e3c", 
    x"5e3e", x"5e40", x"5e43", x"5e45", x"5e47", x"5e49", x"5e4b", x"5e4d", 
    x"5e4f", x"5e51", x"5e54", x"5e56", x"5e58", x"5e5a", x"5e5c", x"5e5e", 
    x"5e60", x"5e62", x"5e64", x"5e67", x"5e69", x"5e6b", x"5e6d", x"5e6f", 
    x"5e71", x"5e73", x"5e75", x"5e78", x"5e7a", x"5e7c", x"5e7e", x"5e80", 
    x"5e82", x"5e84", x"5e86", x"5e89", x"5e8b", x"5e8d", x"5e8f", x"5e91", 
    x"5e93", x"5e95", x"5e97", x"5e99", x"5e9c", x"5e9e", x"5ea0", x"5ea2", 
    x"5ea4", x"5ea6", x"5ea8", x"5eaa", x"5ead", x"5eaf", x"5eb1", x"5eb3", 
    x"5eb5", x"5eb7", x"5eb9", x"5ebb", x"5ebd", x"5ec0", x"5ec2", x"5ec4", 
    x"5ec6", x"5ec8", x"5eca", x"5ecc", x"5ece", x"5ed0", x"5ed3", x"5ed5", 
    x"5ed7", x"5ed9", x"5edb", x"5edd", x"5edf", x"5ee1", x"5ee3", x"5ee6", 
    x"5ee8", x"5eea", x"5eec", x"5eee", x"5ef0", x"5ef2", x"5ef4", x"5ef6", 
    x"5ef8", x"5efb", x"5efd", x"5eff", x"5f01", x"5f03", x"5f05", x"5f07", 
    x"5f09", x"5f0b", x"5f0e", x"5f10", x"5f12", x"5f14", x"5f16", x"5f18", 
    x"5f1a", x"5f1c", x"5f1e", x"5f20", x"5f23", x"5f25", x"5f27", x"5f29", 
    x"5f2b", x"5f2d", x"5f2f", x"5f31", x"5f33", x"5f35", x"5f38", x"5f3a", 
    x"5f3c", x"5f3e", x"5f40", x"5f42", x"5f44", x"5f46", x"5f48", x"5f4a", 
    x"5f4d", x"5f4f", x"5f51", x"5f53", x"5f55", x"5f57", x"5f59", x"5f5b", 
    x"5f5d", x"5f5f", x"5f61", x"5f64", x"5f66", x"5f68", x"5f6a", x"5f6c", 
    x"5f6e", x"5f70", x"5f72", x"5f74", x"5f76", x"5f79", x"5f7b", x"5f7d", 
    x"5f7f", x"5f81", x"5f83", x"5f85", x"5f87", x"5f89", x"5f8b", x"5f8d", 
    x"5f90", x"5f92", x"5f94", x"5f96", x"5f98", x"5f9a", x"5f9c", x"5f9e", 
    x"5fa0", x"5fa2", x"5fa4", x"5fa7", x"5fa9", x"5fab", x"5fad", x"5faf", 
    x"5fb1", x"5fb3", x"5fb5", x"5fb7", x"5fb9", x"5fbb", x"5fbd", x"5fc0", 
    x"5fc2", x"5fc4", x"5fc6", x"5fc8", x"5fca", x"5fcc", x"5fce", x"5fd0", 
    x"5fd2", x"5fd4", x"5fd6", x"5fd9", x"5fdb", x"5fdd", x"5fdf", x"5fe1", 
    x"5fe3", x"5fe5", x"5fe7", x"5fe9", x"5feb", x"5fed", x"5fef", x"5ff2", 
    x"5ff4", x"5ff6", x"5ff8", x"5ffa", x"5ffc", x"5ffe", x"6000", x"6002", 
    x"6004", x"6006", x"6008", x"600a", x"600d", x"600f", x"6011", x"6013", 
    x"6015", x"6017", x"6019", x"601b", x"601d", x"601f", x"6021", x"6023", 
    x"6025", x"6028", x"602a", x"602c", x"602e", x"6030", x"6032", x"6034", 
    x"6036", x"6038", x"603a", x"603c", x"603e", x"6040", x"6042", x"6045", 
    x"6047", x"6049", x"604b", x"604d", x"604f", x"6051", x"6053", x"6055", 
    x"6057", x"6059", x"605b", x"605d", x"605f", x"6061", x"6064", x"6066", 
    x"6068", x"606a", x"606c", x"606e", x"6070", x"6072", x"6074", x"6076", 
    x"6078", x"607a", x"607c", x"607e", x"6080", x"6083", x"6085", x"6087", 
    x"6089", x"608b", x"608d", x"608f", x"6091", x"6093", x"6095", x"6097", 
    x"6099", x"609b", x"609d", x"609f", x"60a1", x"60a4", x"60a6", x"60a8", 
    x"60aa", x"60ac", x"60ae", x"60b0", x"60b2", x"60b4", x"60b6", x"60b8", 
    x"60ba", x"60bc", x"60be", x"60c0", x"60c2", x"60c4", x"60c6", x"60c9", 
    x"60cb", x"60cd", x"60cf", x"60d1", x"60d3", x"60d5", x"60d7", x"60d9", 
    x"60db", x"60dd", x"60df", x"60e1", x"60e3", x"60e5", x"60e7", x"60e9", 
    x"60eb", x"60ee", x"60f0", x"60f2", x"60f4", x"60f6", x"60f8", x"60fa", 
    x"60fc", x"60fe", x"6100", x"6102", x"6104", x"6106", x"6108", x"610a", 
    x"610c", x"610e", x"6110", x"6112", x"6114", x"6117", x"6119", x"611b", 
    x"611d", x"611f", x"6121", x"6123", x"6125", x"6127", x"6129", x"612b", 
    x"612d", x"612f", x"6131", x"6133", x"6135", x"6137", x"6139", x"613b", 
    x"613d", x"613f", x"6141", x"6143", x"6146", x"6148", x"614a", x"614c", 
    x"614e", x"6150", x"6152", x"6154", x"6156", x"6158", x"615a", x"615c", 
    x"615e", x"6160", x"6162", x"6164", x"6166", x"6168", x"616a", x"616c", 
    x"616e", x"6170", x"6172", x"6174", x"6176", x"6179", x"617b", x"617d", 
    x"617f", x"6181", x"6183", x"6185", x"6187", x"6189", x"618b", x"618d", 
    x"618f", x"6191", x"6193", x"6195", x"6197", x"6199", x"619b", x"619d", 
    x"619f", x"61a1", x"61a3", x"61a5", x"61a7", x"61a9", x"61ab", x"61ad", 
    x"61af", x"61b1", x"61b3", x"61b5", x"61b8", x"61ba", x"61bc", x"61be", 
    x"61c0", x"61c2", x"61c4", x"61c6", x"61c8", x"61ca", x"61cc", x"61ce", 
    x"61d0", x"61d2", x"61d4", x"61d6", x"61d8", x"61da", x"61dc", x"61de", 
    x"61e0", x"61e2", x"61e4", x"61e6", x"61e8", x"61ea", x"61ec", x"61ee", 
    x"61f0", x"61f2", x"61f4", x"61f6", x"61f8", x"61fa", x"61fc", x"61fe", 
    x"6200", x"6202", x"6204", x"6206", x"6208", x"620b", x"620d", x"620f", 
    x"6211", x"6213", x"6215", x"6217", x"6219", x"621b", x"621d", x"621f", 
    x"6221", x"6223", x"6225", x"6227", x"6229", x"622b", x"622d", x"622f", 
    x"6231", x"6233", x"6235", x"6237", x"6239", x"623b", x"623d", x"623f", 
    x"6241", x"6243", x"6245", x"6247", x"6249", x"624b", x"624d", x"624f", 
    x"6251", x"6253", x"6255", x"6257", x"6259", x"625b", x"625d", x"625f", 
    x"6261", x"6263", x"6265", x"6267", x"6269", x"626b", x"626d", x"626f", 
    x"6271", x"6273", x"6275", x"6277", x"6279", x"627b", x"627d", x"627f", 
    x"6281", x"6283", x"6285", x"6287", x"6289", x"628b", x"628d", x"628f", 
    x"6291", x"6293", x"6295", x"6297", x"6299", x"629b", x"629d", x"629f", 
    x"62a1", x"62a3", x"62a5", x"62a7", x"62a9", x"62ab", x"62ad", x"62af", 
    x"62b1", x"62b3", x"62b5", x"62b7", x"62b9", x"62bb", x"62bd", x"62bf", 
    x"62c1", x"62c3", x"62c5", x"62c7", x"62c9", x"62cb", x"62cd", x"62cf", 
    x"62d1", x"62d3", x"62d5", x"62d7", x"62d9", x"62db", x"62dd", x"62df", 
    x"62e1", x"62e3", x"62e5", x"62e7", x"62e9", x"62eb", x"62ed", x"62ef", 
    x"62f1", x"62f3", x"62f5", x"62f7", x"62f9", x"62fb", x"62fd", x"62ff", 
    x"6301", x"6303", x"6305", x"6307", x"6309", x"630b", x"630d", x"630f", 
    x"6311", x"6313", x"6315", x"6317", x"6319", x"631b", x"631d", x"631f", 
    x"6321", x"6323", x"6325", x"6327", x"6329", x"632b", x"632d", x"632f", 
    x"6331", x"6333", x"6335", x"6337", x"6339", x"633b", x"633d", x"633f", 
    x"6341", x"6343", x"6345", x"6347", x"6349", x"634b", x"634d", x"634f", 
    x"6351", x"6353", x"6355", x"6357", x"6359", x"635b", x"635d", x"635e", 
    x"6360", x"6362", x"6364", x"6366", x"6368", x"636a", x"636c", x"636e", 
    x"6370", x"6372", x"6374", x"6376", x"6378", x"637a", x"637c", x"637e", 
    x"6380", x"6382", x"6384", x"6386", x"6388", x"638a", x"638c", x"638e", 
    x"6390", x"6392", x"6394", x"6396", x"6398", x"639a", x"639c", x"639e", 
    x"63a0", x"63a2", x"63a4", x"63a6", x"63a8", x"63aa", x"63ac", x"63ae", 
    x"63af", x"63b1", x"63b3", x"63b5", x"63b7", x"63b9", x"63bb", x"63bd", 
    x"63bf", x"63c1", x"63c3", x"63c5", x"63c7", x"63c9", x"63cb", x"63cd", 
    x"63cf", x"63d1", x"63d3", x"63d5", x"63d7", x"63d9", x"63db", x"63dd", 
    x"63df", x"63e1", x"63e3", x"63e5", x"63e7", x"63e9", x"63ea", x"63ec", 
    x"63ee", x"63f0", x"63f2", x"63f4", x"63f6", x"63f8", x"63fa", x"63fc", 
    x"63fe", x"6400", x"6402", x"6404", x"6406", x"6408", x"640a", x"640c", 
    x"640e", x"6410", x"6412", x"6414", x"6416", x"6418", x"641a", x"641c", 
    x"641d", x"641f", x"6421", x"6423", x"6425", x"6427", x"6429", x"642b", 
    x"642d", x"642f", x"6431", x"6433", x"6435", x"6437", x"6439", x"643b", 
    x"643d", x"643f", x"6441", x"6443", x"6445", x"6447", x"6448", x"644a", 
    x"644c", x"644e", x"6450", x"6452", x"6454", x"6456", x"6458", x"645a", 
    x"645c", x"645e", x"6460", x"6462", x"6464", x"6466", x"6468", x"646a", 
    x"646c", x"646e", x"646f", x"6471", x"6473", x"6475", x"6477", x"6479", 
    x"647b", x"647d", x"647f", x"6481", x"6483", x"6485", x"6487", x"6489", 
    x"648b", x"648d", x"648f", x"6491", x"6492", x"6494", x"6496", x"6498", 
    x"649a", x"649c", x"649e", x"64a0", x"64a2", x"64a4", x"64a6", x"64a8", 
    x"64aa", x"64ac", x"64ae", x"64b0", x"64b2", x"64b3", x"64b5", x"64b7", 
    x"64b9", x"64bb", x"64bd", x"64bf", x"64c1", x"64c3", x"64c5", x"64c7", 
    x"64c9", x"64cb", x"64cd", x"64cf", x"64d1", x"64d2", x"64d4", x"64d6", 
    x"64d8", x"64da", x"64dc", x"64de", x"64e0", x"64e2", x"64e4", x"64e6", 
    x"64e8", x"64ea", x"64ec", x"64ee", x"64ef", x"64f1", x"64f3", x"64f5", 
    x"64f7", x"64f9", x"64fb", x"64fd", x"64ff", x"6501", x"6503", x"6505", 
    x"6507", x"6509", x"650a", x"650c", x"650e", x"6510", x"6512", x"6514", 
    x"6516", x"6518", x"651a", x"651c", x"651e", x"6520", x"6522", x"6524", 
    x"6525", x"6527", x"6529", x"652b", x"652d", x"652f", x"6531", x"6533", 
    x"6535", x"6537", x"6539", x"653b", x"653d", x"653e", x"6540", x"6542", 
    x"6544", x"6546", x"6548", x"654a", x"654c", x"654e", x"6550", x"6552", 
    x"6554", x"6556", x"6557", x"6559", x"655b", x"655d", x"655f", x"6561", 
    x"6563", x"6565", x"6567", x"6569", x"656b", x"656d", x"656e", x"6570", 
    x"6572", x"6574", x"6576", x"6578", x"657a", x"657c", x"657e", x"6580", 
    x"6582", x"6584", x"6585", x"6587", x"6589", x"658b", x"658d", x"658f", 
    x"6591", x"6593", x"6595", x"6597", x"6599", x"659a", x"659c", x"659e", 
    x"65a0", x"65a2", x"65a4", x"65a6", x"65a8", x"65aa", x"65ac", x"65ae", 
    x"65af", x"65b1", x"65b3", x"65b5", x"65b7", x"65b9", x"65bb", x"65bd", 
    x"65bf", x"65c1", x"65c3", x"65c4", x"65c6", x"65c8", x"65ca", x"65cc", 
    x"65ce", x"65d0", x"65d2", x"65d4", x"65d6", x"65d7", x"65d9", x"65db", 
    x"65dd", x"65df", x"65e1", x"65e3", x"65e5", x"65e7", x"65e9", x"65ea", 
    x"65ec", x"65ee", x"65f0", x"65f2", x"65f4", x"65f6", x"65f8", x"65fa", 
    x"65fc", x"65fd", x"65ff", x"6601", x"6603", x"6605", x"6607", x"6609", 
    x"660b", x"660d", x"660f", x"6610", x"6612", x"6614", x"6616", x"6618", 
    x"661a", x"661c", x"661e", x"6620", x"6622", x"6623", x"6625", x"6627", 
    x"6629", x"662b", x"662d", x"662f", x"6631", x"6633", x"6634", x"6636", 
    x"6638", x"663a", x"663c", x"663e", x"6640", x"6642", x"6644", x"6645", 
    x"6647", x"6649", x"664b", x"664d", x"664f", x"6651", x"6653", x"6655", 
    x"6656", x"6658", x"665a", x"665c", x"665e", x"6660", x"6662", x"6664", 
    x"6666", x"6667", x"6669", x"666b", x"666d", x"666f", x"6671", x"6673", 
    x"6675", x"6676", x"6678", x"667a", x"667c", x"667e", x"6680", x"6682", 
    x"6684", x"6686", x"6687", x"6689", x"668b", x"668d", x"668f", x"6691", 
    x"6693", x"6695", x"6696", x"6698", x"669a", x"669c", x"669e", x"66a0", 
    x"66a2", x"66a4", x"66a5", x"66a7", x"66a9", x"66ab", x"66ad", x"66af", 
    x"66b1", x"66b3", x"66b4", x"66b6", x"66b8", x"66ba", x"66bc", x"66be", 
    x"66c0", x"66c2", x"66c3", x"66c5", x"66c7", x"66c9", x"66cb", x"66cd", 
    x"66cf", x"66d1", x"66d2", x"66d4", x"66d6", x"66d8", x"66da", x"66dc", 
    x"66de", x"66e0", x"66e1", x"66e3", x"66e5", x"66e7", x"66e9", x"66eb", 
    x"66ed", x"66ee", x"66f0", x"66f2", x"66f4", x"66f6", x"66f8", x"66fa", 
    x"66fc", x"66fd", x"66ff", x"6701", x"6703", x"6705", x"6707", x"6709", 
    x"670a", x"670c", x"670e", x"6710", x"6712", x"6714", x"6716", x"6718", 
    x"6719", x"671b", x"671d", x"671f", x"6721", x"6723", x"6725", x"6726", 
    x"6728", x"672a", x"672c", x"672e", x"6730", x"6732", x"6733", x"6735", 
    x"6737", x"6739", x"673b", x"673d", x"673f", x"6740", x"6742", x"6744", 
    x"6746", x"6748", x"674a", x"674c", x"674d", x"674f", x"6751", x"6753", 
    x"6755", x"6757", x"6759", x"675a", x"675c", x"675e", x"6760", x"6762", 
    x"6764", x"6765", x"6767", x"6769", x"676b", x"676d", x"676f", x"6771", 
    x"6772", x"6774", x"6776", x"6778", x"677a", x"677c", x"677e", x"677f", 
    x"6781", x"6783", x"6785", x"6787", x"6789", x"678a", x"678c", x"678e", 
    x"6790", x"6792", x"6794", x"6796", x"6797", x"6799", x"679b", x"679d", 
    x"679f", x"67a1", x"67a2", x"67a4", x"67a6", x"67a8", x"67aa", x"67ac", 
    x"67ae", x"67af", x"67b1", x"67b3", x"67b5", x"67b7", x"67b9", x"67ba", 
    x"67bc", x"67be", x"67c0", x"67c2", x"67c4", x"67c5", x"67c7", x"67c9", 
    x"67cb", x"67cd", x"67cf", x"67d0", x"67d2", x"67d4", x"67d6", x"67d8", 
    x"67da", x"67dc", x"67dd", x"67df", x"67e1", x"67e3", x"67e5", x"67e7", 
    x"67e8", x"67ea", x"67ec", x"67ee", x"67f0", x"67f2", x"67f3", x"67f5", 
    x"67f7", x"67f9", x"67fb", x"67fd", x"67fe", x"6800", x"6802", x"6804", 
    x"6806", x"6807", x"6809", x"680b", x"680d", x"680f", x"6811", x"6812", 
    x"6814", x"6816", x"6818", x"681a", x"681c", x"681d", x"681f", x"6821", 
    x"6823", x"6825", x"6827", x"6828", x"682a", x"682c", x"682e", x"6830", 
    x"6832", x"6833", x"6835", x"6837", x"6839", x"683b", x"683c", x"683e", 
    x"6840", x"6842", x"6844", x"6846", x"6847", x"6849", x"684b", x"684d", 
    x"684f", x"6851", x"6852", x"6854", x"6856", x"6858", x"685a", x"685b", 
    x"685d", x"685f", x"6861", x"6863", x"6865", x"6866", x"6868", x"686a", 
    x"686c", x"686e", x"686f", x"6871", x"6873", x"6875", x"6877", x"6879", 
    x"687a", x"687c", x"687e", x"6880", x"6882", x"6883", x"6885", x"6887", 
    x"6889", x"688b", x"688c", x"688e", x"6890", x"6892", x"6894", x"6896", 
    x"6897", x"6899", x"689b", x"689d", x"689f", x"68a0", x"68a2", x"68a4", 
    x"68a6", x"68a8", x"68a9", x"68ab", x"68ad", x"68af", x"68b1", x"68b2", 
    x"68b4", x"68b6", x"68b8", x"68ba", x"68bb", x"68bd", x"68bf", x"68c1", 
    x"68c3", x"68c5", x"68c6", x"68c8", x"68ca", x"68cc", x"68ce", x"68cf", 
    x"68d1", x"68d3", x"68d5", x"68d7", x"68d8", x"68da", x"68dc", x"68de", 
    x"68e0", x"68e1", x"68e3", x"68e5", x"68e7", x"68e9", x"68ea", x"68ec", 
    x"68ee", x"68f0", x"68f2", x"68f3", x"68f5", x"68f7", x"68f9", x"68fb", 
    x"68fc", x"68fe", x"6900", x"6902", x"6904", x"6905", x"6907", x"6909", 
    x"690b", x"690d", x"690e", x"6910", x"6912", x"6914", x"6915", x"6917", 
    x"6919", x"691b", x"691d", x"691e", x"6920", x"6922", x"6924", x"6926", 
    x"6927", x"6929", x"692b", x"692d", x"692f", x"6930", x"6932", x"6934", 
    x"6936", x"6938", x"6939", x"693b", x"693d", x"693f", x"6940", x"6942", 
    x"6944", x"6946", x"6948", x"6949", x"694b", x"694d", x"694f", x"6951", 
    x"6952", x"6954", x"6956", x"6958", x"6959", x"695b", x"695d", x"695f", 
    x"6961", x"6962", x"6964", x"6966", x"6968", x"696a", x"696b", x"696d", 
    x"696f", x"6971", x"6972", x"6974", x"6976", x"6978", x"697a", x"697b", 
    x"697d", x"697f", x"6981", x"6982", x"6984", x"6986", x"6988", x"698a", 
    x"698b", x"698d", x"698f", x"6991", x"6992", x"6994", x"6996", x"6998", 
    x"699a", x"699b", x"699d", x"699f", x"69a1", x"69a2", x"69a4", x"69a6", 
    x"69a8", x"69a9", x"69ab", x"69ad", x"69af", x"69b1", x"69b2", x"69b4", 
    x"69b6", x"69b8", x"69b9", x"69bb", x"69bd", x"69bf", x"69c1", x"69c2", 
    x"69c4", x"69c6", x"69c8", x"69c9", x"69cb", x"69cd", x"69cf", x"69d0", 
    x"69d2", x"69d4", x"69d6", x"69d8", x"69d9", x"69db", x"69dd", x"69df", 
    x"69e0", x"69e2", x"69e4", x"69e6", x"69e7", x"69e9", x"69eb", x"69ed", 
    x"69ee", x"69f0", x"69f2", x"69f4", x"69f6", x"69f7", x"69f9", x"69fb", 
    x"69fd", x"69fe", x"6a00", x"6a02", x"6a04", x"6a05", x"6a07", x"6a09", 
    x"6a0b", x"6a0c", x"6a0e", x"6a10", x"6a12", x"6a13", x"6a15", x"6a17", 
    x"6a19", x"6a1a", x"6a1c", x"6a1e", x"6a20", x"6a21", x"6a23", x"6a25", 
    x"6a27", x"6a29", x"6a2a", x"6a2c", x"6a2e", x"6a30", x"6a31", x"6a33", 
    x"6a35", x"6a37", x"6a38", x"6a3a", x"6a3c", x"6a3e", x"6a3f", x"6a41", 
    x"6a43", x"6a45", x"6a46", x"6a48", x"6a4a", x"6a4c", x"6a4d", x"6a4f", 
    x"6a51", x"6a53", x"6a54", x"6a56", x"6a58", x"6a5a", x"6a5b", x"6a5d", 
    x"6a5f", x"6a61", x"6a62", x"6a64", x"6a66", x"6a68", x"6a69", x"6a6b", 
    x"6a6d", x"6a6f", x"6a70", x"6a72", x"6a74", x"6a75", x"6a77", x"6a79", 
    x"6a7b", x"6a7c", x"6a7e", x"6a80", x"6a82", x"6a83", x"6a85", x"6a87", 
    x"6a89", x"6a8a", x"6a8c", x"6a8e", x"6a90", x"6a91", x"6a93", x"6a95", 
    x"6a97", x"6a98", x"6a9a", x"6a9c", x"6a9e", x"6a9f", x"6aa1", x"6aa3", 
    x"6aa4", x"6aa6", x"6aa8", x"6aaa", x"6aab", x"6aad", x"6aaf", x"6ab1", 
    x"6ab2", x"6ab4", x"6ab6", x"6ab8", x"6ab9", x"6abb", x"6abd", x"6abf", 
    x"6ac0", x"6ac2", x"6ac4", x"6ac5", x"6ac7", x"6ac9", x"6acb", x"6acc", 
    x"6ace", x"6ad0", x"6ad2", x"6ad3", x"6ad5", x"6ad7", x"6ad8", x"6ada", 
    x"6adc", x"6ade", x"6adf", x"6ae1", x"6ae3", x"6ae5", x"6ae6", x"6ae8", 
    x"6aea", x"6aec", x"6aed", x"6aef", x"6af1", x"6af2", x"6af4", x"6af6", 
    x"6af8", x"6af9", x"6afb", x"6afd", x"6afe", x"6b00", x"6b02", x"6b04", 
    x"6b05", x"6b07", x"6b09", x"6b0b", x"6b0c", x"6b0e", x"6b10", x"6b11", 
    x"6b13", x"6b15", x"6b17", x"6b18", x"6b1a", x"6b1c", x"6b1d", x"6b1f", 
    x"6b21", x"6b23", x"6b24", x"6b26", x"6b28", x"6b2a", x"6b2b", x"6b2d", 
    x"6b2f", x"6b30", x"6b32", x"6b34", x"6b36", x"6b37", x"6b39", x"6b3b", 
    x"6b3c", x"6b3e", x"6b40", x"6b42", x"6b43", x"6b45", x"6b47", x"6b48", 
    x"6b4a", x"6b4c", x"6b4e", x"6b4f", x"6b51", x"6b53", x"6b54", x"6b56", 
    x"6b58", x"6b5a", x"6b5b", x"6b5d", x"6b5f", x"6b60", x"6b62", x"6b64", 
    x"6b65", x"6b67", x"6b69", x"6b6b", x"6b6c", x"6b6e", x"6b70", x"6b71", 
    x"6b73", x"6b75", x"6b77", x"6b78", x"6b7a", x"6b7c", x"6b7d", x"6b7f", 
    x"6b81", x"6b83", x"6b84", x"6b86", x"6b88", x"6b89", x"6b8b", x"6b8d", 
    x"6b8e", x"6b90", x"6b92", x"6b94", x"6b95", x"6b97", x"6b99", x"6b9a", 
    x"6b9c", x"6b9e", x"6b9f", x"6ba1", x"6ba3", x"6ba5", x"6ba6", x"6ba8", 
    x"6baa", x"6bab", x"6bad", x"6baf", x"6bb0", x"6bb2", x"6bb4", x"6bb6", 
    x"6bb7", x"6bb9", x"6bbb", x"6bbc", x"6bbe", x"6bc0", x"6bc1", x"6bc3", 
    x"6bc5", x"6bc6", x"6bc8", x"6bca", x"6bcc", x"6bcd", x"6bcf", x"6bd1", 
    x"6bd2", x"6bd4", x"6bd6", x"6bd7", x"6bd9", x"6bdb", x"6bdd", x"6bde", 
    x"6be0", x"6be2", x"6be3", x"6be5", x"6be7", x"6be8", x"6bea", x"6bec", 
    x"6bed", x"6bef", x"6bf1", x"6bf2", x"6bf4", x"6bf6", x"6bf8", x"6bf9", 
    x"6bfb", x"6bfd", x"6bfe", x"6c00", x"6c02", x"6c03", x"6c05", x"6c07", 
    x"6c08", x"6c0a", x"6c0c", x"6c0d", x"6c0f", x"6c11", x"6c12", x"6c14", 
    x"6c16", x"6c18", x"6c19", x"6c1b", x"6c1d", x"6c1e", x"6c20", x"6c22", 
    x"6c23", x"6c25", x"6c27", x"6c28", x"6c2a", x"6c2c", x"6c2d", x"6c2f", 
    x"6c31", x"6c32", x"6c34", x"6c36", x"6c37", x"6c39", x"6c3b", x"6c3c", 
    x"6c3e", x"6c40", x"6c42", x"6c43", x"6c45", x"6c47", x"6c48", x"6c4a", 
    x"6c4c", x"6c4d", x"6c4f", x"6c51", x"6c52", x"6c54", x"6c56", x"6c57", 
    x"6c59", x"6c5b", x"6c5c", x"6c5e", x"6c60", x"6c61", x"6c63", x"6c65", 
    x"6c66", x"6c68", x"6c6a", x"6c6b", x"6c6d", x"6c6f", x"6c70", x"6c72", 
    x"6c74", x"6c75", x"6c77", x"6c79", x"6c7a", x"6c7c", x"6c7e", x"6c7f", 
    x"6c81", x"6c83", x"6c84", x"6c86", x"6c88", x"6c89", x"6c8b", x"6c8d", 
    x"6c8e", x"6c90", x"6c92", x"6c93", x"6c95", x"6c97", x"6c98", x"6c9a", 
    x"6c9c", x"6c9d", x"6c9f", x"6ca1", x"6ca2", x"6ca4", x"6ca6", x"6ca7", 
    x"6ca9", x"6cab", x"6cac", x"6cae", x"6cb0", x"6cb1", x"6cb3", x"6cb5", 
    x"6cb6", x"6cb8", x"6cba", x"6cbb", x"6cbd", x"6cbf", x"6cc0", x"6cc2", 
    x"6cc3", x"6cc5", x"6cc7", x"6cc8", x"6cca", x"6ccc", x"6ccd", x"6ccf", 
    x"6cd1", x"6cd2", x"6cd4", x"6cd6", x"6cd7", x"6cd9", x"6cdb", x"6cdc", 
    x"6cde", x"6ce0", x"6ce1", x"6ce3", x"6ce5", x"6ce6", x"6ce8", x"6cea", 
    x"6ceb", x"6ced", x"6cee", x"6cf0", x"6cf2", x"6cf3", x"6cf5", x"6cf7", 
    x"6cf8", x"6cfa", x"6cfc", x"6cfd", x"6cff", x"6d01", x"6d02", x"6d04", 
    x"6d06", x"6d07", x"6d09", x"6d0a", x"6d0c", x"6d0e", x"6d0f", x"6d11", 
    x"6d13", x"6d14", x"6d16", x"6d18", x"6d19", x"6d1b", x"6d1d", x"6d1e", 
    x"6d20", x"6d21", x"6d23", x"6d25", x"6d26", x"6d28", x"6d2a", x"6d2b", 
    x"6d2d", x"6d2f", x"6d30", x"6d32", x"6d34", x"6d35", x"6d37", x"6d38", 
    x"6d3a", x"6d3c", x"6d3d", x"6d3f", x"6d41", x"6d42", x"6d44", x"6d46", 
    x"6d47", x"6d49", x"6d4a", x"6d4c", x"6d4e", x"6d4f", x"6d51", x"6d53", 
    x"6d54", x"6d56", x"6d58", x"6d59", x"6d5b", x"6d5c", x"6d5e", x"6d60", 
    x"6d61", x"6d63", x"6d65", x"6d66", x"6d68", x"6d69", x"6d6b", x"6d6d", 
    x"6d6e", x"6d70", x"6d72", x"6d73", x"6d75", x"6d76", x"6d78", x"6d7a", 
    x"6d7b", x"6d7d", x"6d7f", x"6d80", x"6d82", x"6d84", x"6d85", x"6d87", 
    x"6d88", x"6d8a", x"6d8c", x"6d8d", x"6d8f", x"6d91", x"6d92", x"6d94", 
    x"6d95", x"6d97", x"6d99", x"6d9a", x"6d9c", x"6d9d", x"6d9f", x"6da1", 
    x"6da2", x"6da4", x"6da6", x"6da7", x"6da9", x"6daa", x"6dac", x"6dae", 
    x"6daf", x"6db1", x"6db3", x"6db4", x"6db6", x"6db7", x"6db9", x"6dbb", 
    x"6dbc", x"6dbe", x"6dbf", x"6dc1", x"6dc3", x"6dc4", x"6dc6", x"6dc8", 
    x"6dc9", x"6dcb", x"6dcc", x"6dce", x"6dd0", x"6dd1", x"6dd3", x"6dd4", 
    x"6dd6", x"6dd8", x"6dd9", x"6ddb", x"6ddd", x"6dde", x"6de0", x"6de1", 
    x"6de3", x"6de5", x"6de6", x"6de8", x"6de9", x"6deb", x"6ded", x"6dee", 
    x"6df0", x"6df1", x"6df3", x"6df5", x"6df6", x"6df8", x"6dfa", x"6dfb", 
    x"6dfd", x"6dfe", x"6e00", x"6e02", x"6e03", x"6e05", x"6e06", x"6e08", 
    x"6e0a", x"6e0b", x"6e0d", x"6e0e", x"6e10", x"6e12", x"6e13", x"6e15", 
    x"6e16", x"6e18", x"6e1a", x"6e1b", x"6e1d", x"6e1e", x"6e20", x"6e22", 
    x"6e23", x"6e25", x"6e26", x"6e28", x"6e2a", x"6e2b", x"6e2d", x"6e2e", 
    x"6e30", x"6e32", x"6e33", x"6e35", x"6e36", x"6e38", x"6e3a", x"6e3b", 
    x"6e3d", x"6e3e", x"6e40", x"6e42", x"6e43", x"6e45", x"6e46", x"6e48", 
    x"6e4a", x"6e4b", x"6e4d", x"6e4e", x"6e50", x"6e52", x"6e53", x"6e55", 
    x"6e56", x"6e58", x"6e59", x"6e5b", x"6e5d", x"6e5e", x"6e60", x"6e61", 
    x"6e63", x"6e65", x"6e66", x"6e68", x"6e69", x"6e6b", x"6e6d", x"6e6e", 
    x"6e70", x"6e71", x"6e73", x"6e75", x"6e76", x"6e78", x"6e79", x"6e7b", 
    x"6e7c", x"6e7e", x"6e80", x"6e81", x"6e83", x"6e84", x"6e86", x"6e88", 
    x"6e89", x"6e8b", x"6e8c", x"6e8e", x"6e8f", x"6e91", x"6e93", x"6e94", 
    x"6e96", x"6e97", x"6e99", x"6e9b", x"6e9c", x"6e9e", x"6e9f", x"6ea1", 
    x"6ea2", x"6ea4", x"6ea6", x"6ea7", x"6ea9", x"6eaa", x"6eac", x"6ead", 
    x"6eaf", x"6eb1", x"6eb2", x"6eb4", x"6eb5", x"6eb7", x"6eb9", x"6eba", 
    x"6ebc", x"6ebd", x"6ebf", x"6ec0", x"6ec2", x"6ec4", x"6ec5", x"6ec7", 
    x"6ec8", x"6eca", x"6ecb", x"6ecd", x"6ecf", x"6ed0", x"6ed2", x"6ed3", 
    x"6ed5", x"6ed6", x"6ed8", x"6eda", x"6edb", x"6edd", x"6ede", x"6ee0", 
    x"6ee1", x"6ee3", x"6ee5", x"6ee6", x"6ee8", x"6ee9", x"6eeb", x"6eec", 
    x"6eee", x"6ef0", x"6ef1", x"6ef3", x"6ef4", x"6ef6", x"6ef7", x"6ef9", 
    x"6efb", x"6efc", x"6efe", x"6eff", x"6f01", x"6f02", x"6f04", x"6f05", 
    x"6f07", x"6f09", x"6f0a", x"6f0c", x"6f0d", x"6f0f", x"6f10", x"6f12", 
    x"6f14", x"6f15", x"6f17", x"6f18", x"6f1a", x"6f1b", x"6f1d", x"6f1e", 
    x"6f20", x"6f22", x"6f23", x"6f25", x"6f26", x"6f28", x"6f29", x"6f2b", 
    x"6f2c", x"6f2e", x"6f30", x"6f31", x"6f33", x"6f34", x"6f36", x"6f37", 
    x"6f39", x"6f3a", x"6f3c", x"6f3e", x"6f3f", x"6f41", x"6f42", x"6f44", 
    x"6f45", x"6f47", x"6f48", x"6f4a", x"6f4c", x"6f4d", x"6f4f", x"6f50", 
    x"6f52", x"6f53", x"6f55", x"6f56", x"6f58", x"6f59", x"6f5b", x"6f5d", 
    x"6f5e", x"6f60", x"6f61", x"6f63", x"6f64", x"6f66", x"6f67", x"6f69", 
    x"6f6b", x"6f6c", x"6f6e", x"6f6f", x"6f71", x"6f72", x"6f74", x"6f75", 
    x"6f77", x"6f78", x"6f7a", x"6f7c", x"6f7d", x"6f7f", x"6f80", x"6f82", 
    x"6f83", x"6f85", x"6f86", x"6f88", x"6f89", x"6f8b", x"6f8c", x"6f8e", 
    x"6f90", x"6f91", x"6f93", x"6f94", x"6f96", x"6f97", x"6f99", x"6f9a", 
    x"6f9c", x"6f9d", x"6f9f", x"6fa0", x"6fa2", x"6fa4", x"6fa5", x"6fa7", 
    x"6fa8", x"6faa", x"6fab", x"6fad", x"6fae", x"6fb0", x"6fb1", x"6fb3", 
    x"6fb4", x"6fb6", x"6fb8", x"6fb9", x"6fbb", x"6fbc", x"6fbe", x"6fbf", 
    x"6fc1", x"6fc2", x"6fc4", x"6fc5", x"6fc7", x"6fc8", x"6fca", x"6fcb", 
    x"6fcd", x"6fce", x"6fd0", x"6fd2", x"6fd3", x"6fd5", x"6fd6", x"6fd8", 
    x"6fd9", x"6fdb", x"6fdc", x"6fde", x"6fdf", x"6fe1", x"6fe2", x"6fe4", 
    x"6fe5", x"6fe7", x"6fe8", x"6fea", x"6feb", x"6fed", x"6fef", x"6ff0", 
    x"6ff2", x"6ff3", x"6ff5", x"6ff6", x"6ff8", x"6ff9", x"6ffb", x"6ffc", 
    x"6ffe", x"6fff", x"7001", x"7002", x"7004", x"7005", x"7007", x"7008", 
    x"700a", x"700b", x"700d", x"700e", x"7010", x"7012", x"7013", x"7015", 
    x"7016", x"7018", x"7019", x"701b", x"701c", x"701e", x"701f", x"7021", 
    x"7022", x"7024", x"7025", x"7027", x"7028", x"702a", x"702b", x"702d", 
    x"702e", x"7030", x"7031", x"7033", x"7034", x"7036", x"7037", x"7039", 
    x"703a", x"703c", x"703d", x"703f", x"7040", x"7042", x"7043", x"7045", 
    x"7046", x"7048", x"7049", x"704b", x"704c", x"704e", x"7050", x"7051", 
    x"7053", x"7054", x"7056", x"7057", x"7059", x"705a", x"705c", x"705d", 
    x"705f", x"7060", x"7062", x"7063", x"7065", x"7066", x"7068", x"7069", 
    x"706b", x"706c", x"706e", x"706f", x"7071", x"7072", x"7074", x"7075", 
    x"7077", x"7078", x"707a", x"707b", x"707d", x"707e", x"7080", x"7081", 
    x"7083", x"7084", x"7086", x"7087", x"7089", x"708a", x"708c", x"708d", 
    x"708f", x"7090", x"7092", x"7093", x"7095", x"7096", x"7098", x"7099", 
    x"709b", x"709c", x"709e", x"709f", x"70a0", x"70a2", x"70a3", x"70a5", 
    x"70a6", x"70a8", x"70a9", x"70ab", x"70ac", x"70ae", x"70af", x"70b1", 
    x"70b2", x"70b4", x"70b5", x"70b7", x"70b8", x"70ba", x"70bb", x"70bd", 
    x"70be", x"70c0", x"70c1", x"70c3", x"70c4", x"70c6", x"70c7", x"70c9", 
    x"70ca", x"70cc", x"70cd", x"70cf", x"70d0", x"70d2", x"70d3", x"70d5", 
    x"70d6", x"70d8", x"70d9", x"70db", x"70dc", x"70dd", x"70df", x"70e0", 
    x"70e2", x"70e3", x"70e5", x"70e6", x"70e8", x"70e9", x"70eb", x"70ec", 
    x"70ee", x"70ef", x"70f1", x"70f2", x"70f4", x"70f5", x"70f7", x"70f8", 
    x"70fa", x"70fb", x"70fd", x"70fe", x"70ff", x"7101", x"7102", x"7104", 
    x"7105", x"7107", x"7108", x"710a", x"710b", x"710d", x"710e", x"7110", 
    x"7111", x"7113", x"7114", x"7116", x"7117", x"7119", x"711a", x"711b", 
    x"711d", x"711e", x"7120", x"7121", x"7123", x"7124", x"7126", x"7127", 
    x"7129", x"712a", x"712c", x"712d", x"712f", x"7130", x"7131", x"7133", 
    x"7134", x"7136", x"7137", x"7139", x"713a", x"713c", x"713d", x"713f", 
    x"7140", x"7142", x"7143", x"7145", x"7146", x"7147", x"7149", x"714a", 
    x"714c", x"714d", x"714f", x"7150", x"7152", x"7153", x"7155", x"7156", 
    x"7158", x"7159", x"715a", x"715c", x"715d", x"715f", x"7160", x"7162", 
    x"7163", x"7165", x"7166", x"7168", x"7169", x"716a", x"716c", x"716d", 
    x"716f", x"7170", x"7172", x"7173", x"7175", x"7176", x"7178", x"7179", 
    x"717a", x"717c", x"717d", x"717f", x"7180", x"7182", x"7183", x"7185", 
    x"7186", x"7188", x"7189", x"718a", x"718c", x"718d", x"718f", x"7190", 
    x"7192", x"7193", x"7195", x"7196", x"7197", x"7199", x"719a", x"719c", 
    x"719d", x"719f", x"71a0", x"71a2", x"71a3", x"71a5", x"71a6", x"71a7", 
    x"71a9", x"71aa", x"71ac", x"71ad", x"71af", x"71b0", x"71b2", x"71b3", 
    x"71b4", x"71b6", x"71b7", x"71b9", x"71ba", x"71bc", x"71bd", x"71be", 
    x"71c0", x"71c1", x"71c3", x"71c4", x"71c6", x"71c7", x"71c9", x"71ca", 
    x"71cb", x"71cd", x"71ce", x"71d0", x"71d1", x"71d3", x"71d4", x"71d6", 
    x"71d7", x"71d8", x"71da", x"71db", x"71dd", x"71de", x"71e0", x"71e1", 
    x"71e2", x"71e4", x"71e5", x"71e7", x"71e8", x"71ea", x"71eb", x"71ec", 
    x"71ee", x"71ef", x"71f1", x"71f2", x"71f4", x"71f5", x"71f6", x"71f8", 
    x"71f9", x"71fb", x"71fc", x"71fe", x"71ff", x"7200", x"7202", x"7203", 
    x"7205", x"7206", x"7208", x"7209", x"720a", x"720c", x"720d", x"720f", 
    x"7210", x"7212", x"7213", x"7214", x"7216", x"7217", x"7219", x"721a", 
    x"721c", x"721d", x"721e", x"7220", x"7221", x"7223", x"7224", x"7226", 
    x"7227", x"7228", x"722a", x"722b", x"722d", x"722e", x"722f", x"7231", 
    x"7232", x"7234", x"7235", x"7237", x"7238", x"7239", x"723b", x"723c", 
    x"723e", x"723f", x"7240", x"7242", x"7243", x"7245", x"7246", x"7248", 
    x"7249", x"724a", x"724c", x"724d", x"724f", x"7250", x"7251", x"7253", 
    x"7254", x"7256", x"7257", x"7259", x"725a", x"725b", x"725d", x"725e", 
    x"7260", x"7261", x"7262", x"7264", x"7265", x"7267", x"7268", x"7269", 
    x"726b", x"726c", x"726e", x"726f", x"7270", x"7272", x"7273", x"7275", 
    x"7276", x"7278", x"7279", x"727a", x"727c", x"727d", x"727f", x"7280", 
    x"7281", x"7283", x"7284", x"7286", x"7287", x"7288", x"728a", x"728b", 
    x"728d", x"728e", x"728f", x"7291", x"7292", x"7294", x"7295", x"7296", 
    x"7298", x"7299", x"729b", x"729c", x"729d", x"729f", x"72a0", x"72a2", 
    x"72a3", x"72a4", x"72a6", x"72a7", x"72a9", x"72aa", x"72ab", x"72ad", 
    x"72ae", x"72b0", x"72b1", x"72b2", x"72b4", x"72b5", x"72b6", x"72b8", 
    x"72b9", x"72bb", x"72bc", x"72bd", x"72bf", x"72c0", x"72c2", x"72c3", 
    x"72c4", x"72c6", x"72c7", x"72c9", x"72ca", x"72cb", x"72cd", x"72ce", 
    x"72d0", x"72d1", x"72d2", x"72d4", x"72d5", x"72d6", x"72d8", x"72d9", 
    x"72db", x"72dc", x"72dd", x"72df", x"72e0", x"72e2", x"72e3", x"72e4", 
    x"72e6", x"72e7", x"72e8", x"72ea", x"72eb", x"72ed", x"72ee", x"72ef", 
    x"72f1", x"72f2", x"72f4", x"72f5", x"72f6", x"72f8", x"72f9", x"72fa", 
    x"72fc", x"72fd", x"72ff", x"7300", x"7301", x"7303", x"7304", x"7305", 
    x"7307", x"7308", x"730a", x"730b", x"730c", x"730e", x"730f", x"7311", 
    x"7312", x"7313", x"7315", x"7316", x"7317", x"7319", x"731a", x"731c", 
    x"731d", x"731e", x"7320", x"7321", x"7322", x"7324", x"7325", x"7326", 
    x"7328", x"7329", x"732b", x"732c", x"732d", x"732f", x"7330", x"7331", 
    x"7333", x"7334", x"7336", x"7337", x"7338", x"733a", x"733b", x"733c", 
    x"733e", x"733f", x"7340", x"7342", x"7343", x"7345", x"7346", x"7347", 
    x"7349", x"734a", x"734b", x"734d", x"734e", x"7350", x"7351", x"7352", 
    x"7354", x"7355", x"7356", x"7358", x"7359", x"735a", x"735c", x"735d", 
    x"735e", x"7360", x"7361", x"7363", x"7364", x"7365", x"7367", x"7368", 
    x"7369", x"736b", x"736c", x"736d", x"736f", x"7370", x"7372", x"7373", 
    x"7374", x"7376", x"7377", x"7378", x"737a", x"737b", x"737c", x"737e", 
    x"737f", x"7380", x"7382", x"7383", x"7384", x"7386", x"7387", x"7389", 
    x"738a", x"738b", x"738d", x"738e", x"738f", x"7391", x"7392", x"7393", 
    x"7395", x"7396", x"7397", x"7399", x"739a", x"739b", x"739d", x"739e", 
    x"739f", x"73a1", x"73a2", x"73a4", x"73a5", x"73a6", x"73a8", x"73a9", 
    x"73aa", x"73ac", x"73ad", x"73ae", x"73b0", x"73b1", x"73b2", x"73b4", 
    x"73b5", x"73b6", x"73b8", x"73b9", x"73ba", x"73bc", x"73bd", x"73be", 
    x"73c0", x"73c1", x"73c2", x"73c4", x"73c5", x"73c6", x"73c8", x"73c9", 
    x"73ca", x"73cc", x"73cd", x"73ce", x"73d0", x"73d1", x"73d3", x"73d4", 
    x"73d5", x"73d7", x"73d8", x"73d9", x"73db", x"73dc", x"73dd", x"73df", 
    x"73e0", x"73e1", x"73e3", x"73e4", x"73e5", x"73e7", x"73e8", x"73e9", 
    x"73eb", x"73ec", x"73ed", x"73ef", x"73f0", x"73f1", x"73f3", x"73f4", 
    x"73f5", x"73f7", x"73f8", x"73f9", x"73fa", x"73fc", x"73fd", x"73fe", 
    x"7400", x"7401", x"7402", x"7404", x"7405", x"7406", x"7408", x"7409", 
    x"740a", x"740c", x"740d", x"740e", x"7410", x"7411", x"7412", x"7414", 
    x"7415", x"7416", x"7418", x"7419", x"741a", x"741c", x"741d", x"741e", 
    x"7420", x"7421", x"7422", x"7424", x"7425", x"7426", x"7428", x"7429", 
    x"742a", x"742b", x"742d", x"742e", x"742f", x"7431", x"7432", x"7433", 
    x"7435", x"7436", x"7437", x"7439", x"743a", x"743b", x"743d", x"743e", 
    x"743f", x"7441", x"7442", x"7443", x"7444", x"7446", x"7447", x"7448", 
    x"744a", x"744b", x"744c", x"744e", x"744f", x"7450", x"7452", x"7453", 
    x"7454", x"7456", x"7457", x"7458", x"7459", x"745b", x"745c", x"745d", 
    x"745f", x"7460", x"7461", x"7463", x"7464", x"7465", x"7467", x"7468", 
    x"7469", x"746a", x"746c", x"746d", x"746e", x"7470", x"7471", x"7472", 
    x"7474", x"7475", x"7476", x"7478", x"7479", x"747a", x"747b", x"747d", 
    x"747e", x"747f", x"7481", x"7482", x"7483", x"7485", x"7486", x"7487", 
    x"7488", x"748a", x"748b", x"748c", x"748e", x"748f", x"7490", x"7492", 
    x"7493", x"7494", x"7495", x"7497", x"7498", x"7499", x"749b", x"749c", 
    x"749d", x"749e", x"74a0", x"74a1", x"74a2", x"74a4", x"74a5", x"74a6", 
    x"74a8", x"74a9", x"74aa", x"74ab", x"74ad", x"74ae", x"74af", x"74b1", 
    x"74b2", x"74b3", x"74b4", x"74b6", x"74b7", x"74b8", x"74ba", x"74bb", 
    x"74bc", x"74bd", x"74bf", x"74c0", x"74c1", x"74c3", x"74c4", x"74c5", 
    x"74c6", x"74c8", x"74c9", x"74ca", x"74cc", x"74cd", x"74ce", x"74cf", 
    x"74d1", x"74d2", x"74d3", x"74d5", x"74d6", x"74d7", x"74d8", x"74da", 
    x"74db", x"74dc", x"74de", x"74df", x"74e0", x"74e1", x"74e3", x"74e4", 
    x"74e5", x"74e7", x"74e8", x"74e9", x"74ea", x"74ec", x"74ed", x"74ee", 
    x"74f0", x"74f1", x"74f2", x"74f3", x"74f5", x"74f6", x"74f7", x"74f8", 
    x"74fa", x"74fb", x"74fc", x"74fe", x"74ff", x"7500", x"7501", x"7503", 
    x"7504", x"7505", x"7506", x"7508", x"7509", x"750a", x"750c", x"750d", 
    x"750e", x"750f", x"7511", x"7512", x"7513", x"7514", x"7516", x"7517", 
    x"7518", x"751a", x"751b", x"751c", x"751d", x"751f", x"7520", x"7521", 
    x"7522", x"7524", x"7525", x"7526", x"7527", x"7529", x"752a", x"752b", 
    x"752d", x"752e", x"752f", x"7530", x"7532", x"7533", x"7534", x"7535", 
    x"7537", x"7538", x"7539", x"753a", x"753c", x"753d", x"753e", x"753f", 
    x"7541", x"7542", x"7543", x"7544", x"7546", x"7547", x"7548", x"754a", 
    x"754b", x"754c", x"754d", x"754f", x"7550", x"7551", x"7552", x"7554", 
    x"7555", x"7556", x"7557", x"7559", x"755a", x"755b", x"755c", x"755e", 
    x"755f", x"7560", x"7561", x"7563", x"7564", x"7565", x"7566", x"7568", 
    x"7569", x"756a", x"756b", x"756d", x"756e", x"756f", x"7570", x"7572", 
    x"7573", x"7574", x"7575", x"7577", x"7578", x"7579", x"757a", x"757c", 
    x"757d", x"757e", x"757f", x"7581", x"7582", x"7583", x"7584", x"7586", 
    x"7587", x"7588", x"7589", x"758b", x"758c", x"758d", x"758e", x"7590", 
    x"7591", x"7592", x"7593", x"7594", x"7596", x"7597", x"7598", x"7599", 
    x"759b", x"759c", x"759d", x"759e", x"75a0", x"75a1", x"75a2", x"75a3", 
    x"75a5", x"75a6", x"75a7", x"75a8", x"75aa", x"75ab", x"75ac", x"75ad", 
    x"75ae", x"75b0", x"75b1", x"75b2", x"75b3", x"75b5", x"75b6", x"75b7", 
    x"75b8", x"75ba", x"75bb", x"75bc", x"75bd", x"75bf", x"75c0", x"75c1", 
    x"75c2", x"75c3", x"75c5", x"75c6", x"75c7", x"75c8", x"75ca", x"75cb", 
    x"75cc", x"75cd", x"75cf", x"75d0", x"75d1", x"75d2", x"75d3", x"75d5", 
    x"75d6", x"75d7", x"75d8", x"75da", x"75db", x"75dc", x"75dd", x"75de", 
    x"75e0", x"75e1", x"75e2", x"75e3", x"75e5", x"75e6", x"75e7", x"75e8", 
    x"75e9", x"75eb", x"75ec", x"75ed", x"75ee", x"75f0", x"75f1", x"75f2", 
    x"75f3", x"75f4", x"75f6", x"75f7", x"75f8", x"75f9", x"75fb", x"75fc", 
    x"75fd", x"75fe", x"75ff", x"7601", x"7602", x"7603", x"7604", x"7606", 
    x"7607", x"7608", x"7609", x"760a", x"760c", x"760d", x"760e", x"760f", 
    x"7610", x"7612", x"7613", x"7614", x"7615", x"7617", x"7618", x"7619", 
    x"761a", x"761b", x"761d", x"761e", x"761f", x"7620", x"7621", x"7623", 
    x"7624", x"7625", x"7626", x"7627", x"7629", x"762a", x"762b", x"762c", 
    x"762d", x"762f", x"7630", x"7631", x"7632", x"7634", x"7635", x"7636", 
    x"7637", x"7638", x"763a", x"763b", x"763c", x"763d", x"763e", x"7640", 
    x"7641", x"7642", x"7643", x"7644", x"7646", x"7647", x"7648", x"7649", 
    x"764a", x"764c", x"764d", x"764e", x"764f", x"7650", x"7652", x"7653", 
    x"7654", x"7655", x"7656", x"7658", x"7659", x"765a", x"765b", x"765c", 
    x"765e", x"765f", x"7660", x"7661", x"7662", x"7664", x"7665", x"7666", 
    x"7667", x"7668", x"7669", x"766b", x"766c", x"766d", x"766e", x"766f", 
    x"7671", x"7672", x"7673", x"7674", x"7675", x"7677", x"7678", x"7679", 
    x"767a", x"767b", x"767d", x"767e", x"767f", x"7680", x"7681", x"7682", 
    x"7684", x"7685", x"7686", x"7687", x"7688", x"768a", x"768b", x"768c", 
    x"768d", x"768e", x"768f", x"7691", x"7692", x"7693", x"7694", x"7695", 
    x"7697", x"7698", x"7699", x"769a", x"769b", x"769d", x"769e", x"769f", 
    x"76a0", x"76a1", x"76a2", x"76a4", x"76a5", x"76a6", x"76a7", x"76a8", 
    x"76a9", x"76ab", x"76ac", x"76ad", x"76ae", x"76af", x"76b1", x"76b2", 
    x"76b3", x"76b4", x"76b5", x"76b6", x"76b8", x"76b9", x"76ba", x"76bb", 
    x"76bc", x"76bd", x"76bf", x"76c0", x"76c1", x"76c2", x"76c3", x"76c4", 
    x"76c6", x"76c7", x"76c8", x"76c9", x"76ca", x"76cc", x"76cd", x"76ce", 
    x"76cf", x"76d0", x"76d1", x"76d3", x"76d4", x"76d5", x"76d6", x"76d7", 
    x"76d8", x"76da", x"76db", x"76dc", x"76dd", x"76de", x"76df", x"76e1", 
    x"76e2", x"76e3", x"76e4", x"76e5", x"76e6", x"76e7", x"76e9", x"76ea", 
    x"76eb", x"76ec", x"76ed", x"76ee", x"76f0", x"76f1", x"76f2", x"76f3", 
    x"76f4", x"76f5", x"76f7", x"76f8", x"76f9", x"76fa", x"76fb", x"76fc", 
    x"76fe", x"76ff", x"7700", x"7701", x"7702", x"7703", x"7704", x"7706", 
    x"7707", x"7708", x"7709", x"770a", x"770b", x"770d", x"770e", x"770f", 
    x"7710", x"7711", x"7712", x"7713", x"7715", x"7716", x"7717", x"7718", 
    x"7719", x"771a", x"771c", x"771d", x"771e", x"771f", x"7720", x"7721", 
    x"7722", x"7724", x"7725", x"7726", x"7727", x"7728", x"7729", x"772a", 
    x"772c", x"772d", x"772e", x"772f", x"7730", x"7731", x"7732", x"7734", 
    x"7735", x"7736", x"7737", x"7738", x"7739", x"773a", x"773c", x"773d", 
    x"773e", x"773f", x"7740", x"7741", x"7742", x"7744", x"7745", x"7746", 
    x"7747", x"7748", x"7749", x"774a", x"774c", x"774d", x"774e", x"774f", 
    x"7750", x"7751", x"7752", x"7754", x"7755", x"7756", x"7757", x"7758", 
    x"7759", x"775a", x"775c", x"775d", x"775e", x"775f", x"7760", x"7761", 
    x"7762", x"7763", x"7765", x"7766", x"7767", x"7768", x"7769", x"776a", 
    x"776b", x"776d", x"776e", x"776f", x"7770", x"7771", x"7772", x"7773", 
    x"7774", x"7776", x"7777", x"7778", x"7779", x"777a", x"777b", x"777c", 
    x"777d", x"777f", x"7780", x"7781", x"7782", x"7783", x"7784", x"7785", 
    x"7786", x"7788", x"7789", x"778a", x"778b", x"778c", x"778d", x"778e", 
    x"778f", x"7791", x"7792", x"7793", x"7794", x"7795", x"7796", x"7797", 
    x"7798", x"7799", x"779b", x"779c", x"779d", x"779e", x"779f", x"77a0", 
    x"77a1", x"77a2", x"77a4", x"77a5", x"77a6", x"77a7", x"77a8", x"77a9", 
    x"77aa", x"77ab", x"77ac", x"77ae", x"77af", x"77b0", x"77b1", x"77b2", 
    x"77b3", x"77b4", x"77b5", x"77b6", x"77b8", x"77b9", x"77ba", x"77bb", 
    x"77bc", x"77bd", x"77be", x"77bf", x"77c0", x"77c2", x"77c3", x"77c4", 
    x"77c5", x"77c6", x"77c7", x"77c8", x"77c9", x"77ca", x"77cc", x"77cd", 
    x"77ce", x"77cf", x"77d0", x"77d1", x"77d2", x"77d3", x"77d4", x"77d6", 
    x"77d7", x"77d8", x"77d9", x"77da", x"77db", x"77dc", x"77dd", x"77de", 
    x"77df", x"77e1", x"77e2", x"77e3", x"77e4", x"77e5", x"77e6", x"77e7", 
    x"77e8", x"77e9", x"77ea", x"77ec", x"77ed", x"77ee", x"77ef", x"77f0", 
    x"77f1", x"77f2", x"77f3", x"77f4", x"77f5", x"77f7", x"77f8", x"77f9", 
    x"77fa", x"77fb", x"77fc", x"77fd", x"77fe", x"77ff", x"7800", x"7801", 
    x"7803", x"7804", x"7805", x"7806", x"7807", x"7808", x"7809", x"780a", 
    x"780b", x"780c", x"780d", x"780f", x"7810", x"7811", x"7812", x"7813", 
    x"7814", x"7815", x"7816", x"7817", x"7818", x"7819", x"781a", x"781c", 
    x"781d", x"781e", x"781f", x"7820", x"7821", x"7822", x"7823", x"7824", 
    x"7825", x"7826", x"7828", x"7829", x"782a", x"782b", x"782c", x"782d", 
    x"782e", x"782f", x"7830", x"7831", x"7832", x"7833", x"7834", x"7836", 
    x"7837", x"7838", x"7839", x"783a", x"783b", x"783c", x"783d", x"783e", 
    x"783f", x"7840", x"7841", x"7842", x"7844", x"7845", x"7846", x"7847", 
    x"7848", x"7849", x"784a", x"784b", x"784c", x"784d", x"784e", x"784f", 
    x"7850", x"7852", x"7853", x"7854", x"7855", x"7856", x"7857", x"7858", 
    x"7859", x"785a", x"785b", x"785c", x"785d", x"785e", x"785f", x"7860", 
    x"7862", x"7863", x"7864", x"7865", x"7866", x"7867", x"7868", x"7869", 
    x"786a", x"786b", x"786c", x"786d", x"786e", x"786f", x"7870", x"7872", 
    x"7873", x"7874", x"7875", x"7876", x"7877", x"7878", x"7879", x"787a", 
    x"787b", x"787c", x"787d", x"787e", x"787f", x"7880", x"7881", x"7883", 
    x"7884", x"7885", x"7886", x"7887", x"7888", x"7889", x"788a", x"788b", 
    x"788c", x"788d", x"788e", x"788f", x"7890", x"7891", x"7892", x"7893", 
    x"7894", x"7896", x"7897", x"7898", x"7899", x"789a", x"789b", x"789c", 
    x"789d", x"789e", x"789f", x"78a0", x"78a1", x"78a2", x"78a3", x"78a4", 
    x"78a5", x"78a6", x"78a7", x"78a8", x"78a9", x"78ab", x"78ac", x"78ad", 
    x"78ae", x"78af", x"78b0", x"78b1", x"78b2", x"78b3", x"78b4", x"78b5", 
    x"78b6", x"78b7", x"78b8", x"78b9", x"78ba", x"78bb", x"78bc", x"78bd", 
    x"78be", x"78bf", x"78c0", x"78c2", x"78c3", x"78c4", x"78c5", x"78c6", 
    x"78c7", x"78c8", x"78c9", x"78ca", x"78cb", x"78cc", x"78cd", x"78ce", 
    x"78cf", x"78d0", x"78d1", x"78d2", x"78d3", x"78d4", x"78d5", x"78d6", 
    x"78d7", x"78d8", x"78d9", x"78da", x"78db", x"78dd", x"78de", x"78df", 
    x"78e0", x"78e1", x"78e2", x"78e3", x"78e4", x"78e5", x"78e6", x"78e7", 
    x"78e8", x"78e9", x"78ea", x"78eb", x"78ec", x"78ed", x"78ee", x"78ef", 
    x"78f0", x"78f1", x"78f2", x"78f3", x"78f4", x"78f5", x"78f6", x"78f7", 
    x"78f8", x"78f9", x"78fa", x"78fb", x"78fc", x"78fd", x"78fe", x"7900", 
    x"7901", x"7902", x"7903", x"7904", x"7905", x"7906", x"7907", x"7908", 
    x"7909", x"790a", x"790b", x"790c", x"790d", x"790e", x"790f", x"7910", 
    x"7911", x"7912", x"7913", x"7914", x"7915", x"7916", x"7917", x"7918", 
    x"7919", x"791a", x"791b", x"791c", x"791d", x"791e", x"791f", x"7920", 
    x"7921", x"7922", x"7923", x"7924", x"7925", x"7926", x"7927", x"7928", 
    x"7929", x"792a", x"792b", x"792c", x"792d", x"792e", x"792f", x"7930", 
    x"7931", x"7932", x"7933", x"7934", x"7935", x"7936", x"7937", x"7938", 
    x"7939", x"793a", x"793b", x"793c", x"793d", x"793e", x"793f", x"7940", 
    x"7941", x"7943", x"7944", x"7945", x"7946", x"7947", x"7948", x"7949", 
    x"794a", x"794b", x"794c", x"794d", x"794e", x"794f", x"7950", x"7951", 
    x"7952", x"7953", x"7954", x"7955", x"7956", x"7957", x"7958", x"7959", 
    x"795a", x"795b", x"795c", x"795d", x"795e", x"795f", x"7960", x"7961", 
    x"7962", x"7963", x"7964", x"7965", x"7966", x"7967", x"7968", x"7969", 
    x"796a", x"796b", x"796b", x"796c", x"796d", x"796e", x"796f", x"7970", 
    x"7971", x"7972", x"7973", x"7974", x"7975", x"7976", x"7977", x"7978", 
    x"7979", x"797a", x"797b", x"797c", x"797d", x"797e", x"797f", x"7980", 
    x"7981", x"7982", x"7983", x"7984", x"7985", x"7986", x"7987", x"7988", 
    x"7989", x"798a", x"798b", x"798c", x"798d", x"798e", x"798f", x"7990", 
    x"7991", x"7992", x"7993", x"7994", x"7995", x"7996", x"7997", x"7998", 
    x"7999", x"799a", x"799b", x"799c", x"799d", x"799e", x"799f", x"79a0", 
    x"79a1", x"79a2", x"79a3", x"79a4", x"79a5", x"79a6", x"79a7", x"79a8", 
    x"79a9", x"79aa", x"79ab", x"79ac", x"79ac", x"79ad", x"79ae", x"79af", 
    x"79b0", x"79b1", x"79b2", x"79b3", x"79b4", x"79b5", x"79b6", x"79b7", 
    x"79b8", x"79b9", x"79ba", x"79bb", x"79bc", x"79bd", x"79be", x"79bf", 
    x"79c0", x"79c1", x"79c2", x"79c3", x"79c4", x"79c5", x"79c6", x"79c7", 
    x"79c8", x"79c9", x"79ca", x"79cb", x"79cc", x"79cd", x"79cd", x"79ce", 
    x"79cf", x"79d0", x"79d1", x"79d2", x"79d3", x"79d4", x"79d5", x"79d6", 
    x"79d7", x"79d8", x"79d9", x"79da", x"79db", x"79dc", x"79dd", x"79de", 
    x"79df", x"79e0", x"79e1", x"79e2", x"79e3", x"79e4", x"79e5", x"79e6", 
    x"79e6", x"79e7", x"79e8", x"79e9", x"79ea", x"79eb", x"79ec", x"79ed", 
    x"79ee", x"79ef", x"79f0", x"79f1", x"79f2", x"79f3", x"79f4", x"79f5", 
    x"79f6", x"79f7", x"79f8", x"79f9", x"79fa", x"79fb", x"79fb", x"79fc", 
    x"79fd", x"79fe", x"79ff", x"7a00", x"7a01", x"7a02", x"7a03", x"7a04", 
    x"7a05", x"7a06", x"7a07", x"7a08", x"7a09", x"7a0a", x"7a0b", x"7a0c", 
    x"7a0d", x"7a0e", x"7a0e", x"7a0f", x"7a10", x"7a11", x"7a12", x"7a13", 
    x"7a14", x"7a15", x"7a16", x"7a17", x"7a18", x"7a19", x"7a1a", x"7a1b", 
    x"7a1c", x"7a1d", x"7a1e", x"7a1e", x"7a1f", x"7a20", x"7a21", x"7a22", 
    x"7a23", x"7a24", x"7a25", x"7a26", x"7a27", x"7a28", x"7a29", x"7a2a", 
    x"7a2b", x"7a2c", x"7a2d", x"7a2e", x"7a2e", x"7a2f", x"7a30", x"7a31", 
    x"7a32", x"7a33", x"7a34", x"7a35", x"7a36", x"7a37", x"7a38", x"7a39", 
    x"7a3a", x"7a3b", x"7a3c", x"7a3c", x"7a3d", x"7a3e", x"7a3f", x"7a40", 
    x"7a41", x"7a42", x"7a43", x"7a44", x"7a45", x"7a46", x"7a47", x"7a48", 
    x"7a49", x"7a49", x"7a4a", x"7a4b", x"7a4c", x"7a4d", x"7a4e", x"7a4f", 
    x"7a50", x"7a51", x"7a52", x"7a53", x"7a54", x"7a55", x"7a56", x"7a56", 
    x"7a57", x"7a58", x"7a59", x"7a5a", x"7a5b", x"7a5c", x"7a5d", x"7a5e", 
    x"7a5f", x"7a60", x"7a61", x"7a61", x"7a62", x"7a63", x"7a64", x"7a65", 
    x"7a66", x"7a67", x"7a68", x"7a69", x"7a6a", x"7a6b", x"7a6c", x"7a6d", 
    x"7a6d", x"7a6e", x"7a6f", x"7a70", x"7a71", x"7a72", x"7a73", x"7a74", 
    x"7a75", x"7a76", x"7a77", x"7a78", x"7a78", x"7a79", x"7a7a", x"7a7b", 
    x"7a7c", x"7a7d", x"7a7e", x"7a7f", x"7a80", x"7a81", x"7a82", x"7a82", 
    x"7a83", x"7a84", x"7a85", x"7a86", x"7a87", x"7a88", x"7a89", x"7a8a", 
    x"7a8b", x"7a8c", x"7a8c", x"7a8d", x"7a8e", x"7a8f", x"7a90", x"7a91", 
    x"7a92", x"7a93", x"7a94", x"7a95", x"7a95", x"7a96", x"7a97", x"7a98", 
    x"7a99", x"7a9a", x"7a9b", x"7a9c", x"7a9d", x"7a9e", x"7a9f", x"7a9f", 
    x"7aa0", x"7aa1", x"7aa2", x"7aa3", x"7aa4", x"7aa5", x"7aa6", x"7aa7", 
    x"7aa8", x"7aa8", x"7aa9", x"7aaa", x"7aab", x"7aac", x"7aad", x"7aae", 
    x"7aaf", x"7ab0", x"7ab0", x"7ab1", x"7ab2", x"7ab3", x"7ab4", x"7ab5", 
    x"7ab6", x"7ab7", x"7ab8", x"7ab9", x"7ab9", x"7aba", x"7abb", x"7abc", 
    x"7abd", x"7abe", x"7abf", x"7ac0", x"7ac1", x"7ac1", x"7ac2", x"7ac3", 
    x"7ac4", x"7ac5", x"7ac6", x"7ac7", x"7ac8", x"7ac9", x"7ac9", x"7aca", 
    x"7acb", x"7acc", x"7acd", x"7ace", x"7acf", x"7ad0", x"7ad1", x"7ad1", 
    x"7ad2", x"7ad3", x"7ad4", x"7ad5", x"7ad6", x"7ad7", x"7ad8", x"7ad8", 
    x"7ad9", x"7ada", x"7adb", x"7adc", x"7add", x"7ade", x"7adf", x"7ae0", 
    x"7ae0", x"7ae1", x"7ae2", x"7ae3", x"7ae4", x"7ae5", x"7ae6", x"7ae7", 
    x"7ae7", x"7ae8", x"7ae9", x"7aea", x"7aeb", x"7aec", x"7aed", x"7aee", 
    x"7aee", x"7aef", x"7af0", x"7af1", x"7af2", x"7af3", x"7af4", x"7af5", 
    x"7af5", x"7af6", x"7af7", x"7af8", x"7af9", x"7afa", x"7afb", x"7afc", 
    x"7afc", x"7afd", x"7afe", x"7aff", x"7b00", x"7b01", x"7b02", x"7b02", 
    x"7b03", x"7b04", x"7b05", x"7b06", x"7b07", x"7b08", x"7b09", x"7b09", 
    x"7b0a", x"7b0b", x"7b0c", x"7b0d", x"7b0e", x"7b0f", x"7b0f", x"7b10", 
    x"7b11", x"7b12", x"7b13", x"7b14", x"7b15", x"7b16", x"7b16", x"7b17", 
    x"7b18", x"7b19", x"7b1a", x"7b1b", x"7b1c", x"7b1c", x"7b1d", x"7b1e", 
    x"7b1f", x"7b20", x"7b21", x"7b22", x"7b22", x"7b23", x"7b24", x"7b25", 
    x"7b26", x"7b27", x"7b28", x"7b28", x"7b29", x"7b2a", x"7b2b", x"7b2c", 
    x"7b2d", x"7b2e", x"7b2e", x"7b2f", x"7b30", x"7b31", x"7b32", x"7b33", 
    x"7b33", x"7b34", x"7b35", x"7b36", x"7b37", x"7b38", x"7b39", x"7b39", 
    x"7b3a", x"7b3b", x"7b3c", x"7b3d", x"7b3e", x"7b3f", x"7b3f", x"7b40", 
    x"7b41", x"7b42", x"7b43", x"7b44", x"7b44", x"7b45", x"7b46", x"7b47", 
    x"7b48", x"7b49", x"7b4a", x"7b4a", x"7b4b", x"7b4c", x"7b4d", x"7b4e", 
    x"7b4f", x"7b4f", x"7b50", x"7b51", x"7b52", x"7b53", x"7b54", x"7b54", 
    x"7b55", x"7b56", x"7b57", x"7b58", x"7b59", x"7b5a", x"7b5a", x"7b5b", 
    x"7b5c", x"7b5d", x"7b5e", x"7b5f", x"7b5f", x"7b60", x"7b61", x"7b62", 
    x"7b63", x"7b64", x"7b64", x"7b65", x"7b66", x"7b67", x"7b68", x"7b69", 
    x"7b69", x"7b6a", x"7b6b", x"7b6c", x"7b6d", x"7b6e", x"7b6e", x"7b6f", 
    x"7b70", x"7b71", x"7b72", x"7b73", x"7b73", x"7b74", x"7b75", x"7b76", 
    x"7b77", x"7b78", x"7b78", x"7b79", x"7b7a", x"7b7b", x"7b7c", x"7b7d", 
    x"7b7d", x"7b7e", x"7b7f", x"7b80", x"7b81", x"7b81", x"7b82", x"7b83", 
    x"7b84", x"7b85", x"7b86", x"7b86", x"7b87", x"7b88", x"7b89", x"7b8a", 
    x"7b8b", x"7b8b", x"7b8c", x"7b8d", x"7b8e", x"7b8f", x"7b8f", x"7b90", 
    x"7b91", x"7b92", x"7b93", x"7b94", x"7b94", x"7b95", x"7b96", x"7b97", 
    x"7b98", x"7b98", x"7b99", x"7b9a", x"7b9b", x"7b9c", x"7b9d", x"7b9d", 
    x"7b9e", x"7b9f", x"7ba0", x"7ba1", x"7ba1", x"7ba2", x"7ba3", x"7ba4", 
    x"7ba5", x"7ba5", x"7ba6", x"7ba7", x"7ba8", x"7ba9", x"7baa", x"7baa", 
    x"7bab", x"7bac", x"7bad", x"7bae", x"7bae", x"7baf", x"7bb0", x"7bb1", 
    x"7bb2", x"7bb2", x"7bb3", x"7bb4", x"7bb5", x"7bb6", x"7bb6", x"7bb7", 
    x"7bb8", x"7bb9", x"7bba", x"7bba", x"7bbb", x"7bbc", x"7bbd", x"7bbe", 
    x"7bbf", x"7bbf", x"7bc0", x"7bc1", x"7bc2", x"7bc3", x"7bc3", x"7bc4", 
    x"7bc5", x"7bc6", x"7bc7", x"7bc7", x"7bc8", x"7bc9", x"7bca", x"7bcb", 
    x"7bcb", x"7bcc", x"7bcd", x"7bce", x"7bcf", x"7bcf", x"7bd0", x"7bd1", 
    x"7bd2", x"7bd2", x"7bd3", x"7bd4", x"7bd5", x"7bd6", x"7bd6", x"7bd7", 
    x"7bd8", x"7bd9", x"7bda", x"7bda", x"7bdb", x"7bdc", x"7bdd", x"7bde", 
    x"7bde", x"7bdf", x"7be0", x"7be1", x"7be2", x"7be2", x"7be3", x"7be4", 
    x"7be5", x"7be6", x"7be6", x"7be7", x"7be8", x"7be9", x"7be9", x"7bea", 
    x"7beb", x"7bec", x"7bed", x"7bed", x"7bee", x"7bef", x"7bf0", x"7bf1", 
    x"7bf1", x"7bf2", x"7bf3", x"7bf4", x"7bf4", x"7bf5", x"7bf6", x"7bf7", 
    x"7bf8", x"7bf8", x"7bf9", x"7bfa", x"7bfb", x"7bfb", x"7bfc", x"7bfd", 
    x"7bfe", x"7bff", x"7bff", x"7c00", x"7c01", x"7c02", x"7c02", x"7c03", 
    x"7c04", x"7c05", x"7c06", x"7c06", x"7c07", x"7c08", x"7c09", x"7c09", 
    x"7c0a", x"7c0b", x"7c0c", x"7c0d", x"7c0d", x"7c0e", x"7c0f", x"7c10", 
    x"7c10", x"7c11", x"7c12", x"7c13", x"7c14", x"7c14", x"7c15", x"7c16", 
    x"7c17", x"7c17", x"7c18", x"7c19", x"7c1a", x"7c1a", x"7c1b", x"7c1c", 
    x"7c1d", x"7c1e", x"7c1e", x"7c1f", x"7c20", x"7c21", x"7c21", x"7c22", 
    x"7c23", x"7c24", x"7c24", x"7c25", x"7c26", x"7c27", x"7c27", x"7c28", 
    x"7c29", x"7c2a", x"7c2b", x"7c2b", x"7c2c", x"7c2d", x"7c2e", x"7c2e", 
    x"7c2f", x"7c30", x"7c31", x"7c31", x"7c32", x"7c33", x"7c34", x"7c34", 
    x"7c35", x"7c36", x"7c37", x"7c37", x"7c38", x"7c39", x"7c3a", x"7c3a", 
    x"7c3b", x"7c3c", x"7c3d", x"7c3e", x"7c3e", x"7c3f", x"7c40", x"7c41", 
    x"7c41", x"7c42", x"7c43", x"7c44", x"7c44", x"7c45", x"7c46", x"7c47", 
    x"7c47", x"7c48", x"7c49", x"7c4a", x"7c4a", x"7c4b", x"7c4c", x"7c4d", 
    x"7c4d", x"7c4e", x"7c4f", x"7c50", x"7c50", x"7c51", x"7c52", x"7c53", 
    x"7c53", x"7c54", x"7c55", x"7c56", x"7c56", x"7c57", x"7c58", x"7c59", 
    x"7c59", x"7c5a", x"7c5b", x"7c5c", x"7c5c", x"7c5d", x"7c5e", x"7c5e", 
    x"7c5f", x"7c60", x"7c61", x"7c61", x"7c62", x"7c63", x"7c64", x"7c64", 
    x"7c65", x"7c66", x"7c67", x"7c67", x"7c68", x"7c69", x"7c6a", x"7c6a", 
    x"7c6b", x"7c6c", x"7c6d", x"7c6d", x"7c6e", x"7c6f", x"7c6f", x"7c70", 
    x"7c71", x"7c72", x"7c72", x"7c73", x"7c74", x"7c75", x"7c75", x"7c76", 
    x"7c77", x"7c78", x"7c78", x"7c79", x"7c7a", x"7c7a", x"7c7b", x"7c7c", 
    x"7c7d", x"7c7d", x"7c7e", x"7c7f", x"7c80", x"7c80", x"7c81", x"7c82", 
    x"7c83", x"7c83", x"7c84", x"7c85", x"7c85", x"7c86", x"7c87", x"7c88", 
    x"7c88", x"7c89", x"7c8a", x"7c8a", x"7c8b", x"7c8c", x"7c8d", x"7c8d", 
    x"7c8e", x"7c8f", x"7c90", x"7c90", x"7c91", x"7c92", x"7c92", x"7c93", 
    x"7c94", x"7c95", x"7c95", x"7c96", x"7c97", x"7c98", x"7c98", x"7c99", 
    x"7c9a", x"7c9a", x"7c9b", x"7c9c", x"7c9d", x"7c9d", x"7c9e", x"7c9f", 
    x"7c9f", x"7ca0", x"7ca1", x"7ca2", x"7ca2", x"7ca3", x"7ca4", x"7ca4", 
    x"7ca5", x"7ca6", x"7ca7", x"7ca7", x"7ca8", x"7ca9", x"7ca9", x"7caa", 
    x"7cab", x"7cac", x"7cac", x"7cad", x"7cae", x"7cae", x"7caf", x"7cb0", 
    x"7cb1", x"7cb1", x"7cb2", x"7cb3", x"7cb3", x"7cb4", x"7cb5", x"7cb5", 
    x"7cb6", x"7cb7", x"7cb8", x"7cb8", x"7cb9", x"7cba", x"7cba", x"7cbb", 
    x"7cbc", x"7cbd", x"7cbd", x"7cbe", x"7cbf", x"7cbf", x"7cc0", x"7cc1", 
    x"7cc1", x"7cc2", x"7cc3", x"7cc4", x"7cc4", x"7cc5", x"7cc6", x"7cc6", 
    x"7cc7", x"7cc8", x"7cc8", x"7cc9", x"7cca", x"7ccb", x"7ccb", x"7ccc", 
    x"7ccd", x"7ccd", x"7cce", x"7ccf", x"7ccf", x"7cd0", x"7cd1", x"7cd2", 
    x"7cd2", x"7cd3", x"7cd4", x"7cd4", x"7cd5", x"7cd6", x"7cd6", x"7cd7", 
    x"7cd8", x"7cd8", x"7cd9", x"7cda", x"7cdb", x"7cdb", x"7cdc", x"7cdd", 
    x"7cdd", x"7cde", x"7cdf", x"7cdf", x"7ce0", x"7ce1", x"7ce1", x"7ce2", 
    x"7ce3", x"7ce4", x"7ce4", x"7ce5", x"7ce6", x"7ce6", x"7ce7", x"7ce8", 
    x"7ce8", x"7ce9", x"7cea", x"7cea", x"7ceb", x"7cec", x"7cec", x"7ced", 
    x"7cee", x"7cee", x"7cef", x"7cf0", x"7cf1", x"7cf1", x"7cf2", x"7cf3", 
    x"7cf3", x"7cf4", x"7cf5", x"7cf5", x"7cf6", x"7cf7", x"7cf7", x"7cf8", 
    x"7cf9", x"7cf9", x"7cfa", x"7cfb", x"7cfb", x"7cfc", x"7cfd", x"7cfd", 
    x"7cfe", x"7cff", x"7cff", x"7d00", x"7d01", x"7d02", x"7d02", x"7d03", 
    x"7d04", x"7d04", x"7d05", x"7d06", x"7d06", x"7d07", x"7d08", x"7d08", 
    x"7d09", x"7d0a", x"7d0a", x"7d0b", x"7d0c", x"7d0c", x"7d0d", x"7d0e", 
    x"7d0e", x"7d0f", x"7d10", x"7d10", x"7d11", x"7d12", x"7d12", x"7d13", 
    x"7d14", x"7d14", x"7d15", x"7d16", x"7d16", x"7d17", x"7d18", x"7d18", 
    x"7d19", x"7d1a", x"7d1a", x"7d1b", x"7d1c", x"7d1c", x"7d1d", x"7d1e", 
    x"7d1e", x"7d1f", x"7d20", x"7d20", x"7d21", x"7d22", x"7d22", x"7d23", 
    x"7d24", x"7d24", x"7d25", x"7d26", x"7d26", x"7d27", x"7d28", x"7d28", 
    x"7d29", x"7d29", x"7d2a", x"7d2b", x"7d2b", x"7d2c", x"7d2d", x"7d2d", 
    x"7d2e", x"7d2f", x"7d2f", x"7d30", x"7d31", x"7d31", x"7d32", x"7d33", 
    x"7d33", x"7d34", x"7d35", x"7d35", x"7d36", x"7d37", x"7d37", x"7d38", 
    x"7d39", x"7d39", x"7d3a", x"7d3a", x"7d3b", x"7d3c", x"7d3c", x"7d3d", 
    x"7d3e", x"7d3e", x"7d3f", x"7d40", x"7d40", x"7d41", x"7d42", x"7d42", 
    x"7d43", x"7d44", x"7d44", x"7d45", x"7d45", x"7d46", x"7d47", x"7d47", 
    x"7d48", x"7d49", x"7d49", x"7d4a", x"7d4b", x"7d4b", x"7d4c", x"7d4d", 
    x"7d4d", x"7d4e", x"7d4e", x"7d4f", x"7d50", x"7d50", x"7d51", x"7d52", 
    x"7d52", x"7d53", x"7d54", x"7d54", x"7d55", x"7d56", x"7d56", x"7d57", 
    x"7d57", x"7d58", x"7d59", x"7d59", x"7d5a", x"7d5b", x"7d5b", x"7d5c", 
    x"7d5c", x"7d5d", x"7d5e", x"7d5e", x"7d5f", x"7d60", x"7d60", x"7d61", 
    x"7d62", x"7d62", x"7d63", x"7d63", x"7d64", x"7d65", x"7d65", x"7d66", 
    x"7d67", x"7d67", x"7d68", x"7d68", x"7d69", x"7d6a", x"7d6a", x"7d6b", 
    x"7d6c", x"7d6c", x"7d6d", x"7d6e", x"7d6e", x"7d6f", x"7d6f", x"7d70", 
    x"7d71", x"7d71", x"7d72", x"7d73", x"7d73", x"7d74", x"7d74", x"7d75", 
    x"7d76", x"7d76", x"7d77", x"7d77", x"7d78", x"7d79", x"7d79", x"7d7a", 
    x"7d7b", x"7d7b", x"7d7c", x"7d7c", x"7d7d", x"7d7e", x"7d7e", x"7d7f", 
    x"7d80", x"7d80", x"7d81", x"7d81", x"7d82", x"7d83", x"7d83", x"7d84", 
    x"7d84", x"7d85", x"7d86", x"7d86", x"7d87", x"7d88", x"7d88", x"7d89", 
    x"7d89", x"7d8a", x"7d8b", x"7d8b", x"7d8c", x"7d8c", x"7d8d", x"7d8e", 
    x"7d8e", x"7d8f", x"7d90", x"7d90", x"7d91", x"7d91", x"7d92", x"7d93", 
    x"7d93", x"7d94", x"7d94", x"7d95", x"7d96", x"7d96", x"7d97", x"7d97", 
    x"7d98", x"7d99", x"7d99", x"7d9a", x"7d9a", x"7d9b", x"7d9c", x"7d9c", 
    x"7d9d", x"7d9d", x"7d9e", x"7d9f", x"7d9f", x"7da0", x"7da0", x"7da1", 
    x"7da2", x"7da2", x"7da3", x"7da3", x"7da4", x"7da5", x"7da5", x"7da6", 
    x"7da6", x"7da7", x"7da8", x"7da8", x"7da9", x"7da9", x"7daa", x"7dab", 
    x"7dab", x"7dac", x"7dac", x"7dad", x"7dae", x"7dae", x"7daf", x"7daf", 
    x"7db0", x"7db1", x"7db1", x"7db2", x"7db2", x"7db3", x"7db4", x"7db4", 
    x"7db5", x"7db5", x"7db6", x"7db7", x"7db7", x"7db8", x"7db8", x"7db9", 
    x"7db9", x"7dba", x"7dbb", x"7dbb", x"7dbc", x"7dbc", x"7dbd", x"7dbe", 
    x"7dbe", x"7dbf", x"7dbf", x"7dc0", x"7dc1", x"7dc1", x"7dc2", x"7dc2", 
    x"7dc3", x"7dc3", x"7dc4", x"7dc5", x"7dc5", x"7dc6", x"7dc6", x"7dc7", 
    x"7dc8", x"7dc8", x"7dc9", x"7dc9", x"7dca", x"7dca", x"7dcb", x"7dcc", 
    x"7dcc", x"7dcd", x"7dcd", x"7dce", x"7dce", x"7dcf", x"7dd0", x"7dd0", 
    x"7dd1", x"7dd1", x"7dd2", x"7dd3", x"7dd3", x"7dd4", x"7dd4", x"7dd5", 
    x"7dd5", x"7dd6", x"7dd7", x"7dd7", x"7dd8", x"7dd8", x"7dd9", x"7dd9", 
    x"7dda", x"7ddb", x"7ddb", x"7ddc", x"7ddc", x"7ddd", x"7ddd", x"7dde", 
    x"7ddf", x"7ddf", x"7de0", x"7de0", x"7de1", x"7de1", x"7de2", x"7de3", 
    x"7de3", x"7de4", x"7de4", x"7de5", x"7de5", x"7de6", x"7de7", x"7de7", 
    x"7de8", x"7de8", x"7de9", x"7de9", x"7dea", x"7dea", x"7deb", x"7dec", 
    x"7dec", x"7ded", x"7ded", x"7dee", x"7dee", x"7def", x"7df0", x"7df0", 
    x"7df1", x"7df1", x"7df2", x"7df2", x"7df3", x"7df3", x"7df4", x"7df5", 
    x"7df5", x"7df6", x"7df6", x"7df7", x"7df7", x"7df8", x"7df8", x"7df9", 
    x"7dfa", x"7dfa", x"7dfb", x"7dfb", x"7dfc", x"7dfc", x"7dfd", x"7dfd", 
    x"7dfe", x"7dff", x"7dff", x"7e00", x"7e00", x"7e01", x"7e01", x"7e02", 
    x"7e02", x"7e03", x"7e04", x"7e04", x"7e05", x"7e05", x"7e06", x"7e06", 
    x"7e07", x"7e07", x"7e08", x"7e09", x"7e09", x"7e0a", x"7e0a", x"7e0b", 
    x"7e0b", x"7e0c", x"7e0c", x"7e0d", x"7e0d", x"7e0e", x"7e0f", x"7e0f", 
    x"7e10", x"7e10", x"7e11", x"7e11", x"7e12", x"7e12", x"7e13", x"7e13", 
    x"7e14", x"7e15", x"7e15", x"7e16", x"7e16", x"7e17", x"7e17", x"7e18", 
    x"7e18", x"7e19", x"7e19", x"7e1a", x"7e1a", x"7e1b", x"7e1c", x"7e1c", 
    x"7e1d", x"7e1d", x"7e1e", x"7e1e", x"7e1f", x"7e1f", x"7e20", x"7e20", 
    x"7e21", x"7e21", x"7e22", x"7e22", x"7e23", x"7e24", x"7e24", x"7e25", 
    x"7e25", x"7e26", x"7e26", x"7e27", x"7e27", x"7e28", x"7e28", x"7e29", 
    x"7e29", x"7e2a", x"7e2a", x"7e2b", x"7e2c", x"7e2c", x"7e2d", x"7e2d", 
    x"7e2e", x"7e2e", x"7e2f", x"7e2f", x"7e30", x"7e30", x"7e31", x"7e31", 
    x"7e32", x"7e32", x"7e33", x"7e33", x"7e34", x"7e34", x"7e35", x"7e36", 
    x"7e36", x"7e37", x"7e37", x"7e38", x"7e38", x"7e39", x"7e39", x"7e3a", 
    x"7e3a", x"7e3b", x"7e3b", x"7e3c", x"7e3c", x"7e3d", x"7e3d", x"7e3e", 
    x"7e3e", x"7e3f", x"7e3f", x"7e40", x"7e40", x"7e41", x"7e41", x"7e42", 
    x"7e42", x"7e43", x"7e44", x"7e44", x"7e45", x"7e45", x"7e46", x"7e46", 
    x"7e47", x"7e47", x"7e48", x"7e48", x"7e49", x"7e49", x"7e4a", x"7e4a", 
    x"7e4b", x"7e4b", x"7e4c", x"7e4c", x"7e4d", x"7e4d", x"7e4e", x"7e4e", 
    x"7e4f", x"7e4f", x"7e50", x"7e50", x"7e51", x"7e51", x"7e52", x"7e52", 
    x"7e53", x"7e53", x"7e54", x"7e54", x"7e55", x"7e55", x"7e56", x"7e56", 
    x"7e57", x"7e57", x"7e58", x"7e58", x"7e59", x"7e59", x"7e5a", x"7e5a", 
    x"7e5b", x"7e5b", x"7e5c", x"7e5c", x"7e5d", x"7e5d", x"7e5e", x"7e5e", 
    x"7e5f", x"7e5f", x"7e60", x"7e60", x"7e61", x"7e61", x"7e62", x"7e62", 
    x"7e63", x"7e63", x"7e64", x"7e64", x"7e65", x"7e65", x"7e66", x"7e66", 
    x"7e67", x"7e67", x"7e68", x"7e68", x"7e69", x"7e69", x"7e6a", x"7e6a", 
    x"7e6b", x"7e6b", x"7e6c", x"7e6c", x"7e6d", x"7e6d", x"7e6e", x"7e6e", 
    x"7e6f", x"7e6f", x"7e70", x"7e70", x"7e71", x"7e71", x"7e72", x"7e72", 
    x"7e73", x"7e73", x"7e74", x"7e74", x"7e75", x"7e75", x"7e76", x"7e76", 
    x"7e77", x"7e77", x"7e77", x"7e78", x"7e78", x"7e79", x"7e79", x"7e7a", 
    x"7e7a", x"7e7b", x"7e7b", x"7e7c", x"7e7c", x"7e7d", x"7e7d", x"7e7e", 
    x"7e7e", x"7e7f", x"7e7f", x"7e80", x"7e80", x"7e81", x"7e81", x"7e82", 
    x"7e82", x"7e83", x"7e83", x"7e83", x"7e84", x"7e84", x"7e85", x"7e85", 
    x"7e86", x"7e86", x"7e87", x"7e87", x"7e88", x"7e88", x"7e89", x"7e89", 
    x"7e8a", x"7e8a", x"7e8b", x"7e8b", x"7e8c", x"7e8c", x"7e8d", x"7e8d", 
    x"7e8d", x"7e8e", x"7e8e", x"7e8f", x"7e8f", x"7e90", x"7e90", x"7e91", 
    x"7e91", x"7e92", x"7e92", x"7e93", x"7e93", x"7e94", x"7e94", x"7e94", 
    x"7e95", x"7e95", x"7e96", x"7e96", x"7e97", x"7e97", x"7e98", x"7e98", 
    x"7e99", x"7e99", x"7e9a", x"7e9a", x"7e9b", x"7e9b", x"7e9b", x"7e9c", 
    x"7e9c", x"7e9d", x"7e9d", x"7e9e", x"7e9e", x"7e9f", x"7e9f", x"7ea0", 
    x"7ea0", x"7ea0", x"7ea1", x"7ea1", x"7ea2", x"7ea2", x"7ea3", x"7ea3", 
    x"7ea4", x"7ea4", x"7ea5", x"7ea5", x"7ea6", x"7ea6", x"7ea6", x"7ea7", 
    x"7ea7", x"7ea8", x"7ea8", x"7ea9", x"7ea9", x"7eaa", x"7eaa", x"7eaa", 
    x"7eab", x"7eab", x"7eac", x"7eac", x"7ead", x"7ead", x"7eae", x"7eae", 
    x"7eaf", x"7eaf", x"7eaf", x"7eb0", x"7eb0", x"7eb1", x"7eb1", x"7eb2", 
    x"7eb2", x"7eb3", x"7eb3", x"7eb3", x"7eb4", x"7eb4", x"7eb5", x"7eb5", 
    x"7eb6", x"7eb6", x"7eb7", x"7eb7", x"7eb7", x"7eb8", x"7eb8", x"7eb9", 
    x"7eb9", x"7eba", x"7eba", x"7ebb", x"7ebb", x"7ebb", x"7ebc", x"7ebc", 
    x"7ebd", x"7ebd", x"7ebe", x"7ebe", x"7ebf", x"7ebf", x"7ebf", x"7ec0", 
    x"7ec0", x"7ec1", x"7ec1", x"7ec2", x"7ec2", x"7ec2", x"7ec3", x"7ec3", 
    x"7ec4", x"7ec4", x"7ec5", x"7ec5", x"7ec5", x"7ec6", x"7ec6", x"7ec7", 
    x"7ec7", x"7ec8", x"7ec8", x"7ec9", x"7ec9", x"7ec9", x"7eca", x"7eca", 
    x"7ecb", x"7ecb", x"7ecc", x"7ecc", x"7ecc", x"7ecd", x"7ecd", x"7ece", 
    x"7ece", x"7ecf", x"7ecf", x"7ecf", x"7ed0", x"7ed0", x"7ed1", x"7ed1", 
    x"7ed2", x"7ed2", x"7ed2", x"7ed3", x"7ed3", x"7ed4", x"7ed4", x"7ed4", 
    x"7ed5", x"7ed5", x"7ed6", x"7ed6", x"7ed7", x"7ed7", x"7ed7", x"7ed8", 
    x"7ed8", x"7ed9", x"7ed9", x"7eda", x"7eda", x"7eda", x"7edb", x"7edb", 
    x"7edc", x"7edc", x"7edc", x"7edd", x"7edd", x"7ede", x"7ede", x"7edf", 
    x"7edf", x"7edf", x"7ee0", x"7ee0", x"7ee1", x"7ee1", x"7ee1", x"7ee2", 
    x"7ee2", x"7ee3", x"7ee3", x"7ee4", x"7ee4", x"7ee4", x"7ee5", x"7ee5", 
    x"7ee6", x"7ee6", x"7ee6", x"7ee7", x"7ee7", x"7ee8", x"7ee8", x"7ee8", 
    x"7ee9", x"7ee9", x"7eea", x"7eea", x"7eea", x"7eeb", x"7eeb", x"7eec", 
    x"7eec", x"7eed", x"7eed", x"7eed", x"7eee", x"7eee", x"7eef", x"7eef", 
    x"7eef", x"7ef0", x"7ef0", x"7ef1", x"7ef1", x"7ef1", x"7ef2", x"7ef2", 
    x"7ef3", x"7ef3", x"7ef3", x"7ef4", x"7ef4", x"7ef5", x"7ef5", x"7ef5", 
    x"7ef6", x"7ef6", x"7ef7", x"7ef7", x"7ef7", x"7ef8", x"7ef8", x"7ef9", 
    x"7ef9", x"7ef9", x"7efa", x"7efa", x"7efb", x"7efb", x"7efb", x"7efc", 
    x"7efc", x"7efd", x"7efd", x"7efd", x"7efe", x"7efe", x"7efe", x"7eff", 
    x"7eff", x"7f00", x"7f00", x"7f00", x"7f01", x"7f01", x"7f02", x"7f02", 
    x"7f02", x"7f03", x"7f03", x"7f04", x"7f04", x"7f04", x"7f05", x"7f05", 
    x"7f05", x"7f06", x"7f06", x"7f07", x"7f07", x"7f07", x"7f08", x"7f08", 
    x"7f09", x"7f09", x"7f09", x"7f0a", x"7f0a", x"7f0a", x"7f0b", x"7f0b", 
    x"7f0c", x"7f0c", x"7f0c", x"7f0d", x"7f0d", x"7f0e", x"7f0e", x"7f0e", 
    x"7f0f", x"7f0f", x"7f0f", x"7f10", x"7f10", x"7f11", x"7f11", x"7f11", 
    x"7f12", x"7f12", x"7f12", x"7f13", x"7f13", x"7f14", x"7f14", x"7f14", 
    x"7f15", x"7f15", x"7f15", x"7f16", x"7f16", x"7f17", x"7f17", x"7f17", 
    x"7f18", x"7f18", x"7f18", x"7f19", x"7f19", x"7f1a", x"7f1a", x"7f1a", 
    x"7f1b", x"7f1b", x"7f1b", x"7f1c", x"7f1c", x"7f1d", x"7f1d", x"7f1d", 
    x"7f1e", x"7f1e", x"7f1e", x"7f1f", x"7f1f", x"7f1f", x"7f20", x"7f20", 
    x"7f21", x"7f21", x"7f21", x"7f22", x"7f22", x"7f22", x"7f23", x"7f23", 
    x"7f23", x"7f24", x"7f24", x"7f25", x"7f25", x"7f25", x"7f26", x"7f26", 
    x"7f26", x"7f27", x"7f27", x"7f27", x"7f28", x"7f28", x"7f29", x"7f29", 
    x"7f29", x"7f2a", x"7f2a", x"7f2a", x"7f2b", x"7f2b", x"7f2b", x"7f2c", 
    x"7f2c", x"7f2c", x"7f2d", x"7f2d", x"7f2e", x"7f2e", x"7f2e", x"7f2f", 
    x"7f2f", x"7f2f", x"7f30", x"7f30", x"7f30", x"7f31", x"7f31", x"7f31", 
    x"7f32", x"7f32", x"7f32", x"7f33", x"7f33", x"7f34", x"7f34", x"7f34", 
    x"7f35", x"7f35", x"7f35", x"7f36", x"7f36", x"7f36", x"7f37", x"7f37", 
    x"7f37", x"7f38", x"7f38", x"7f38", x"7f39", x"7f39", x"7f39", x"7f3a", 
    x"7f3a", x"7f3a", x"7f3b", x"7f3b", x"7f3b", x"7f3c", x"7f3c", x"7f3d", 
    x"7f3d", x"7f3d", x"7f3e", x"7f3e", x"7f3e", x"7f3f", x"7f3f", x"7f3f", 
    x"7f40", x"7f40", x"7f40", x"7f41", x"7f41", x"7f41", x"7f42", x"7f42", 
    x"7f42", x"7f43", x"7f43", x"7f43", x"7f44", x"7f44", x"7f44", x"7f45", 
    x"7f45", x"7f45", x"7f46", x"7f46", x"7f46", x"7f47", x"7f47", x"7f47", 
    x"7f48", x"7f48", x"7f48", x"7f49", x"7f49", x"7f49", x"7f4a", x"7f4a", 
    x"7f4a", x"7f4b", x"7f4b", x"7f4b", x"7f4c", x"7f4c", x"7f4c", x"7f4d", 
    x"7f4d", x"7f4d", x"7f4e", x"7f4e", x"7f4e", x"7f4f", x"7f4f", x"7f4f", 
    x"7f50", x"7f50", x"7f50", x"7f50", x"7f51", x"7f51", x"7f51", x"7f52", 
    x"7f52", x"7f52", x"7f53", x"7f53", x"7f53", x"7f54", x"7f54", x"7f54", 
    x"7f55", x"7f55", x"7f55", x"7f56", x"7f56", x"7f56", x"7f57", x"7f57", 
    x"7f57", x"7f58", x"7f58", x"7f58", x"7f58", x"7f59", x"7f59", x"7f59", 
    x"7f5a", x"7f5a", x"7f5a", x"7f5b", x"7f5b", x"7f5b", x"7f5c", x"7f5c", 
    x"7f5c", x"7f5d", x"7f5d", x"7f5d", x"7f5e", x"7f5e", x"7f5e", x"7f5e", 
    x"7f5f", x"7f5f", x"7f5f", x"7f60", x"7f60", x"7f60", x"7f61", x"7f61", 
    x"7f61", x"7f62", x"7f62", x"7f62", x"7f62", x"7f63", x"7f63", x"7f63", 
    x"7f64", x"7f64", x"7f64", x"7f65", x"7f65", x"7f65", x"7f65", x"7f66", 
    x"7f66", x"7f66", x"7f67", x"7f67", x"7f67", x"7f68", x"7f68", x"7f68", 
    x"7f69", x"7f69", x"7f69", x"7f69", x"7f6a", x"7f6a", x"7f6a", x"7f6b", 
    x"7f6b", x"7f6b", x"7f6c", x"7f6c", x"7f6c", x"7f6c", x"7f6d", x"7f6d", 
    x"7f6d", x"7f6e", x"7f6e", x"7f6e", x"7f6e", x"7f6f", x"7f6f", x"7f6f", 
    x"7f70", x"7f70", x"7f70", x"7f71", x"7f71", x"7f71", x"7f71", x"7f72", 
    x"7f72", x"7f72", x"7f73", x"7f73", x"7f73", x"7f73", x"7f74", x"7f74", 
    x"7f74", x"7f75", x"7f75", x"7f75", x"7f75", x"7f76", x"7f76", x"7f76", 
    x"7f77", x"7f77", x"7f77", x"7f77", x"7f78", x"7f78", x"7f78", x"7f79", 
    x"7f79", x"7f79", x"7f79", x"7f7a", x"7f7a", x"7f7a", x"7f7b", x"7f7b", 
    x"7f7b", x"7f7b", x"7f7c", x"7f7c", x"7f7c", x"7f7d", x"7f7d", x"7f7d", 
    x"7f7d", x"7f7e", x"7f7e", x"7f7e", x"7f7f", x"7f7f", x"7f7f", x"7f7f", 
    x"7f80", x"7f80", x"7f80", x"7f80", x"7f81", x"7f81", x"7f81", x"7f82", 
    x"7f82", x"7f82", x"7f82", x"7f83", x"7f83", x"7f83", x"7f83", x"7f84", 
    x"7f84", x"7f84", x"7f85", x"7f85", x"7f85", x"7f85", x"7f86", x"7f86", 
    x"7f86", x"7f86", x"7f87", x"7f87", x"7f87", x"7f88", x"7f88", x"7f88", 
    x"7f88", x"7f89", x"7f89", x"7f89", x"7f89", x"7f8a", x"7f8a", x"7f8a", 
    x"7f8a", x"7f8b", x"7f8b", x"7f8b", x"7f8c", x"7f8c", x"7f8c", x"7f8c", 
    x"7f8d", x"7f8d", x"7f8d", x"7f8d", x"7f8e", x"7f8e", x"7f8e", x"7f8e", 
    x"7f8f", x"7f8f", x"7f8f", x"7f8f", x"7f90", x"7f90", x"7f90", x"7f90", 
    x"7f91", x"7f91", x"7f91", x"7f91", x"7f92", x"7f92", x"7f92", x"7f93", 
    x"7f93", x"7f93", x"7f93", x"7f94", x"7f94", x"7f94", x"7f94", x"7f95", 
    x"7f95", x"7f95", x"7f95", x"7f96", x"7f96", x"7f96", x"7f96", x"7f97", 
    x"7f97", x"7f97", x"7f97", x"7f98", x"7f98", x"7f98", x"7f98", x"7f99", 
    x"7f99", x"7f99", x"7f99", x"7f9a", x"7f9a", x"7f9a", x"7f9a", x"7f9b", 
    x"7f9b", x"7f9b", x"7f9b", x"7f9c", x"7f9c", x"7f9c", x"7f9c", x"7f9c", 
    x"7f9d", x"7f9d", x"7f9d", x"7f9d", x"7f9e", x"7f9e", x"7f9e", x"7f9e", 
    x"7f9f", x"7f9f", x"7f9f", x"7f9f", x"7fa0", x"7fa0", x"7fa0", x"7fa0", 
    x"7fa1", x"7fa1", x"7fa1", x"7fa1", x"7fa2", x"7fa2", x"7fa2", x"7fa2", 
    x"7fa2", x"7fa3", x"7fa3", x"7fa3", x"7fa3", x"7fa4", x"7fa4", x"7fa4", 
    x"7fa4", x"7fa5", x"7fa5", x"7fa5", x"7fa5", x"7fa6", x"7fa6", x"7fa6", 
    x"7fa6", x"7fa6", x"7fa7", x"7fa7", x"7fa7", x"7fa7", x"7fa8", x"7fa8", 
    x"7fa8", x"7fa8", x"7fa9", x"7fa9", x"7fa9", x"7fa9", x"7fa9", x"7faa", 
    x"7faa", x"7faa", x"7faa", x"7fab", x"7fab", x"7fab", x"7fab", x"7fab", 
    x"7fac", x"7fac", x"7fac", x"7fac", x"7fad", x"7fad", x"7fad", x"7fad", 
    x"7fad", x"7fae", x"7fae", x"7fae", x"7fae", x"7faf", x"7faf", x"7faf", 
    x"7faf", x"7faf", x"7fb0", x"7fb0", x"7fb0", x"7fb0", x"7fb1", x"7fb1", 
    x"7fb1", x"7fb1", x"7fb1", x"7fb2", x"7fb2", x"7fb2", x"7fb2", x"7fb2", 
    x"7fb3", x"7fb3", x"7fb3", x"7fb3", x"7fb4", x"7fb4", x"7fb4", x"7fb4", 
    x"7fb4", x"7fb5", x"7fb5", x"7fb5", x"7fb5", x"7fb5", x"7fb6", x"7fb6", 
    x"7fb6", x"7fb6", x"7fb6", x"7fb7", x"7fb7", x"7fb7", x"7fb7", x"7fb8", 
    x"7fb8", x"7fb8", x"7fb8", x"7fb8", x"7fb9", x"7fb9", x"7fb9", x"7fb9", 
    x"7fb9", x"7fba", x"7fba", x"7fba", x"7fba", x"7fba", x"7fbb", x"7fbb", 
    x"7fbb", x"7fbb", x"7fbb", x"7fbc", x"7fbc", x"7fbc", x"7fbc", x"7fbc", 
    x"7fbd", x"7fbd", x"7fbd", x"7fbd", x"7fbd", x"7fbe", x"7fbe", x"7fbe", 
    x"7fbe", x"7fbe", x"7fbf", x"7fbf", x"7fbf", x"7fbf", x"7fbf", x"7fc0", 
    x"7fc0", x"7fc0", x"7fc0", x"7fc0", x"7fc1", x"7fc1", x"7fc1", x"7fc1", 
    x"7fc1", x"7fc2", x"7fc2", x"7fc2", x"7fc2", x"7fc2", x"7fc2", x"7fc3", 
    x"7fc3", x"7fc3", x"7fc3", x"7fc3", x"7fc4", x"7fc4", x"7fc4", x"7fc4", 
    x"7fc4", x"7fc5", x"7fc5", x"7fc5", x"7fc5", x"7fc5", x"7fc6", x"7fc6", 
    x"7fc6", x"7fc6", x"7fc6", x"7fc6", x"7fc7", x"7fc7", x"7fc7", x"7fc7", 
    x"7fc7", x"7fc8", x"7fc8", x"7fc8", x"7fc8", x"7fc8", x"7fc8", x"7fc9", 
    x"7fc9", x"7fc9", x"7fc9", x"7fc9", x"7fca", x"7fca", x"7fca", x"7fca", 
    x"7fca", x"7fca", x"7fcb", x"7fcb", x"7fcb", x"7fcb", x"7fcb", x"7fcb", 
    x"7fcc", x"7fcc", x"7fcc", x"7fcc", x"7fcc", x"7fcd", x"7fcd", x"7fcd", 
    x"7fcd", x"7fcd", x"7fcd", x"7fce", x"7fce", x"7fce", x"7fce", x"7fce", 
    x"7fce", x"7fcf", x"7fcf", x"7fcf", x"7fcf", x"7fcf", x"7fcf", x"7fd0", 
    x"7fd0", x"7fd0", x"7fd0", x"7fd0", x"7fd0", x"7fd1", x"7fd1", x"7fd1", 
    x"7fd1", x"7fd1", x"7fd1", x"7fd2", x"7fd2", x"7fd2", x"7fd2", x"7fd2", 
    x"7fd2", x"7fd3", x"7fd3", x"7fd3", x"7fd3", x"7fd3", x"7fd3", x"7fd4", 
    x"7fd4", x"7fd4", x"7fd4", x"7fd4", x"7fd4", x"7fd5", x"7fd5", x"7fd5", 
    x"7fd5", x"7fd5", x"7fd5", x"7fd6", x"7fd6", x"7fd6", x"7fd6", x"7fd6", 
    x"7fd6", x"7fd6", x"7fd7", x"7fd7", x"7fd7", x"7fd7", x"7fd7", x"7fd7", 
    x"7fd8", x"7fd8", x"7fd8", x"7fd8", x"7fd8", x"7fd8", x"7fd8", x"7fd9", 
    x"7fd9", x"7fd9", x"7fd9", x"7fd9", x"7fd9", x"7fda", x"7fda", x"7fda", 
    x"7fda", x"7fda", x"7fda", x"7fda", x"7fdb", x"7fdb", x"7fdb", x"7fdb", 
    x"7fdb", x"7fdb", x"7fdb", x"7fdc", x"7fdc", x"7fdc", x"7fdc", x"7fdc", 
    x"7fdc", x"7fdc", x"7fdd", x"7fdd", x"7fdd", x"7fdd", x"7fdd", x"7fdd", 
    x"7fdd", x"7fde", x"7fde", x"7fde", x"7fde", x"7fde", x"7fde", x"7fde", 
    x"7fdf", x"7fdf", x"7fdf", x"7fdf", x"7fdf", x"7fdf", x"7fdf", x"7fe0", 
    x"7fe0", x"7fe0", x"7fe0", x"7fe0", x"7fe0", x"7fe0", x"7fe1", x"7fe1", 
    x"7fe1", x"7fe1", x"7fe1", x"7fe1", x"7fe1", x"7fe1", x"7fe2", x"7fe2", 
    x"7fe2", x"7fe2", x"7fe2", x"7fe2", x"7fe2", x"7fe3", x"7fe3", x"7fe3", 
    x"7fe3", x"7fe3", x"7fe3", x"7fe3", x"7fe3", x"7fe4", x"7fe4", x"7fe4", 
    x"7fe4", x"7fe4", x"7fe4", x"7fe4", x"7fe4", x"7fe5", x"7fe5", x"7fe5", 
    x"7fe5", x"7fe5", x"7fe5", x"7fe5", x"7fe5", x"7fe6", x"7fe6", x"7fe6", 
    x"7fe6", x"7fe6", x"7fe6", x"7fe6", x"7fe6", x"7fe7", x"7fe7", x"7fe7", 
    x"7fe7", x"7fe7", x"7fe7", x"7fe7", x"7fe7", x"7fe8", x"7fe8", x"7fe8", 
    x"7fe8", x"7fe8", x"7fe8", x"7fe8", x"7fe8", x"7fe8", x"7fe9", x"7fe9", 
    x"7fe9", x"7fe9", x"7fe9", x"7fe9", x"7fe9", x"7fe9", x"7fe9", x"7fea", 
    x"7fea", x"7fea", x"7fea", x"7fea", x"7fea", x"7fea", x"7fea", x"7fea", 
    x"7feb", x"7feb", x"7feb", x"7feb", x"7feb", x"7feb", x"7feb", x"7feb", 
    x"7feb", x"7fec", x"7fec", x"7fec", x"7fec", x"7fec", x"7fec", x"7fec", 
    x"7fec", x"7fec", x"7fed", x"7fed", x"7fed", x"7fed", x"7fed", x"7fed", 
    x"7fed", x"7fed", x"7fed", x"7fed", x"7fee", x"7fee", x"7fee", x"7fee", 
    x"7fee", x"7fee", x"7fee", x"7fee", x"7fee", x"7fef", x"7fef", x"7fef", 
    x"7fef", x"7fef", x"7fef", x"7fef", x"7fef", x"7fef", x"7fef", x"7fef", 
    x"7ff0", x"7ff0", x"7ff0", x"7ff0", x"7ff0", x"7ff0", x"7ff0", x"7ff0", 
    x"7ff0", x"7ff0", x"7ff1", x"7ff1", x"7ff1", x"7ff1", x"7ff1", x"7ff1", 
    x"7ff1", x"7ff1", x"7ff1", x"7ff1", x"7ff1", x"7ff2", x"7ff2", x"7ff2", 
    x"7ff2", x"7ff2", x"7ff2", x"7ff2", x"7ff2", x"7ff2", x"7ff2", x"7ff2", 
    x"7ff3", x"7ff3", x"7ff3", x"7ff3", x"7ff3", x"7ff3", x"7ff3", x"7ff3", 
    x"7ff3", x"7ff3", x"7ff3", x"7ff3", x"7ff4", x"7ff4", x"7ff4", x"7ff4", 
    x"7ff4", x"7ff4", x"7ff4", x"7ff4", x"7ff4", x"7ff4", x"7ff4", x"7ff4", 
    x"7ff5", x"7ff5", x"7ff5", x"7ff5", x"7ff5", x"7ff5", x"7ff5", x"7ff5", 
    x"7ff5", x"7ff5", x"7ff5", x"7ff5", x"7ff5", x"7ff6", x"7ff6", x"7ff6", 
    x"7ff6", x"7ff6", x"7ff6", x"7ff6", x"7ff6", x"7ff6", x"7ff6", x"7ff6", 
    x"7ff6", x"7ff6", x"7ff6", x"7ff7", x"7ff7", x"7ff7", x"7ff7", x"7ff7", 
    x"7ff7", x"7ff7", x"7ff7", x"7ff7", x"7ff7", x"7ff7", x"7ff7", x"7ff7", 
    x"7ff7", x"7ff8", x"7ff8", x"7ff8", x"7ff8", x"7ff8", x"7ff8", x"7ff8", 
    x"7ff8", x"7ff8", x"7ff8", x"7ff8", x"7ff8", x"7ff8", x"7ff8", x"7ff8", 
    x"7ff8", x"7ff9", x"7ff9", x"7ff9", x"7ff9", x"7ff9", x"7ff9", x"7ff9", 
    x"7ff9", x"7ff9", x"7ff9", x"7ff9", x"7ff9", x"7ff9", x"7ff9", x"7ff9", 
    x"7ff9", x"7ffa", x"7ffa", x"7ffa", x"7ffa", x"7ffa", x"7ffa", x"7ffa", 
    x"7ffa", x"7ffa", x"7ffa", x"7ffa", x"7ffa", x"7ffa", x"7ffa", x"7ffa", 
    x"7ffa", x"7ffa", x"7ffa", x"7ffa", x"7ffb", x"7ffb", x"7ffb", x"7ffb", 
    x"7ffb", x"7ffb", x"7ffb", x"7ffb", x"7ffb", x"7ffb", x"7ffb", x"7ffb", 
    x"7ffb", x"7ffb", x"7ffb", x"7ffb", x"7ffb", x"7ffb", x"7ffb", x"7ffb", 
    x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", 
    x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", 
    x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", 
    x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", 
    x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", 
    x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", 
    x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffe", x"7ffe", x"7ffe", 
    x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", 
    x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", 
    x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", 
    x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", 
    x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7fff", 
    x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", 
    x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", 
    x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", 
    x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", 
    x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", 
    x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", 
    x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", 
    x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", 
    x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", 
    x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", 
    x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", 
    x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", 
    x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", 
    x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", 
    x"7fff", x"7fff", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", 
    x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", 
    x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", 
    x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", 
    x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", 
    x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffd", x"7ffd", x"7ffd", x"7ffd", 
    x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", 
    x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", 
    x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", 
    x"7ffd", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", 
    x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", 
    x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", 
    x"7ffc", x"7ffb", x"7ffb", x"7ffb", x"7ffb", x"7ffb", x"7ffb", x"7ffb", 
    x"7ffb", x"7ffb", x"7ffb", x"7ffb", x"7ffb", x"7ffb", x"7ffb", x"7ffb", 
    x"7ffb", x"7ffb", x"7ffb", x"7ffb", x"7ffb", x"7ffa", x"7ffa", x"7ffa", 
    x"7ffa", x"7ffa", x"7ffa", x"7ffa", x"7ffa", x"7ffa", x"7ffa", x"7ffa", 
    x"7ffa", x"7ffa", x"7ffa", x"7ffa", x"7ffa", x"7ffa", x"7ffa", x"7ffa", 
    x"7ff9", x"7ff9", x"7ff9", x"7ff9", x"7ff9", x"7ff9", x"7ff9", x"7ff9", 
    x"7ff9", x"7ff9", x"7ff9", x"7ff9", x"7ff9", x"7ff9", x"7ff9", x"7ff9", 
    x"7ff8", x"7ff8", x"7ff8", x"7ff8", x"7ff8", x"7ff8", x"7ff8", x"7ff8", 
    x"7ff8", x"7ff8", x"7ff8", x"7ff8", x"7ff8", x"7ff8", x"7ff8", x"7ff8", 
    x"7ff7", x"7ff7", x"7ff7", x"7ff7", x"7ff7", x"7ff7", x"7ff7", x"7ff7", 
    x"7ff7", x"7ff7", x"7ff7", x"7ff7", x"7ff7", x"7ff7", x"7ff6", x"7ff6", 
    x"7ff6", x"7ff6", x"7ff6", x"7ff6", x"7ff6", x"7ff6", x"7ff6", x"7ff6", 
    x"7ff6", x"7ff6", x"7ff6", x"7ff6", x"7ff5", x"7ff5", x"7ff5", x"7ff5", 
    x"7ff5", x"7ff5", x"7ff5", x"7ff5", x"7ff5", x"7ff5", x"7ff5", x"7ff5", 
    x"7ff5", x"7ff4", x"7ff4", x"7ff4", x"7ff4", x"7ff4", x"7ff4", x"7ff4", 
    x"7ff4", x"7ff4", x"7ff4", x"7ff4", x"7ff4", x"7ff3", x"7ff3", x"7ff3", 
    x"7ff3", x"7ff3", x"7ff3", x"7ff3", x"7ff3", x"7ff3", x"7ff3", x"7ff3", 
    x"7ff3", x"7ff2", x"7ff2", x"7ff2", x"7ff2", x"7ff2", x"7ff2", x"7ff2", 
    x"7ff2", x"7ff2", x"7ff2", x"7ff2", x"7ff1", x"7ff1", x"7ff1", x"7ff1", 
    x"7ff1", x"7ff1", x"7ff1", x"7ff1", x"7ff1", x"7ff1", x"7ff1", x"7ff0", 
    x"7ff0", x"7ff0", x"7ff0", x"7ff0", x"7ff0", x"7ff0", x"7ff0", x"7ff0", 
    x"7ff0", x"7fef", x"7fef", x"7fef", x"7fef", x"7fef", x"7fef", x"7fef", 
    x"7fef", x"7fef", x"7fef", x"7fef", x"7fee", x"7fee", x"7fee", x"7fee", 
    x"7fee", x"7fee", x"7fee", x"7fee", x"7fee", x"7fed", x"7fed", x"7fed", 
    x"7fed", x"7fed", x"7fed", x"7fed", x"7fed", x"7fed", x"7fed", x"7fec", 
    x"7fec", x"7fec", x"7fec", x"7fec", x"7fec", x"7fec", x"7fec", x"7fec", 
    x"7feb", x"7feb", x"7feb", x"7feb", x"7feb", x"7feb", x"7feb", x"7feb", 
    x"7feb", x"7fea", x"7fea", x"7fea", x"7fea", x"7fea", x"7fea", x"7fea", 
    x"7fea", x"7fea", x"7fe9", x"7fe9", x"7fe9", x"7fe9", x"7fe9", x"7fe9", 
    x"7fe9", x"7fe9", x"7fe9", x"7fe8", x"7fe8", x"7fe8", x"7fe8", x"7fe8", 
    x"7fe8", x"7fe8", x"7fe8", x"7fe8", x"7fe7", x"7fe7", x"7fe7", x"7fe7", 
    x"7fe7", x"7fe7", x"7fe7", x"7fe7", x"7fe6", x"7fe6", x"7fe6", x"7fe6", 
    x"7fe6", x"7fe6", x"7fe6", x"7fe6", x"7fe5", x"7fe5", x"7fe5", x"7fe5", 
    x"7fe5", x"7fe5", x"7fe5", x"7fe5", x"7fe4", x"7fe4", x"7fe4", x"7fe4", 
    x"7fe4", x"7fe4", x"7fe4", x"7fe4", x"7fe3", x"7fe3", x"7fe3", x"7fe3", 
    x"7fe3", x"7fe3", x"7fe3", x"7fe3", x"7fe2", x"7fe2", x"7fe2", x"7fe2", 
    x"7fe2", x"7fe2", x"7fe2", x"7fe1", x"7fe1", x"7fe1", x"7fe1", x"7fe1", 
    x"7fe1", x"7fe1", x"7fe1", x"7fe0", x"7fe0", x"7fe0", x"7fe0", x"7fe0", 
    x"7fe0", x"7fe0", x"7fdf", x"7fdf", x"7fdf", x"7fdf", x"7fdf", x"7fdf", 
    x"7fdf", x"7fde", x"7fde", x"7fde", x"7fde", x"7fde", x"7fde", x"7fde", 
    x"7fdd", x"7fdd", x"7fdd", x"7fdd", x"7fdd", x"7fdd", x"7fdd", x"7fdc", 
    x"7fdc", x"7fdc", x"7fdc", x"7fdc", x"7fdc", x"7fdc", x"7fdb", x"7fdb", 
    x"7fdb", x"7fdb", x"7fdb", x"7fdb", x"7fdb", x"7fda", x"7fda", x"7fda", 
    x"7fda", x"7fda", x"7fda", x"7fda", x"7fd9", x"7fd9", x"7fd9", x"7fd9", 
    x"7fd9", x"7fd9", x"7fd8", x"7fd8", x"7fd8", x"7fd8", x"7fd8", x"7fd8", 
    x"7fd8", x"7fd7", x"7fd7", x"7fd7", x"7fd7", x"7fd7", x"7fd7", x"7fd6", 
    x"7fd6", x"7fd6", x"7fd6", x"7fd6", x"7fd6", x"7fd6", x"7fd5", x"7fd5", 
    x"7fd5", x"7fd5", x"7fd5", x"7fd5", x"7fd4", x"7fd4", x"7fd4", x"7fd4", 
    x"7fd4", x"7fd4", x"7fd3", x"7fd3", x"7fd3", x"7fd3", x"7fd3", x"7fd3", 
    x"7fd2", x"7fd2", x"7fd2", x"7fd2", x"7fd2", x"7fd2", x"7fd1", x"7fd1", 
    x"7fd1", x"7fd1", x"7fd1", x"7fd1", x"7fd0", x"7fd0", x"7fd0", x"7fd0", 
    x"7fd0", x"7fd0", x"7fcf", x"7fcf", x"7fcf", x"7fcf", x"7fcf", x"7fcf", 
    x"7fce", x"7fce", x"7fce", x"7fce", x"7fce", x"7fce", x"7fcd", x"7fcd", 
    x"7fcd", x"7fcd", x"7fcd", x"7fcd", x"7fcc", x"7fcc", x"7fcc", x"7fcc", 
    x"7fcc", x"7fcb", x"7fcb", x"7fcb", x"7fcb", x"7fcb", x"7fcb", x"7fca", 
    x"7fca", x"7fca", x"7fca", x"7fca", x"7fca", x"7fc9", x"7fc9", x"7fc9", 
    x"7fc9", x"7fc9", x"7fc8", x"7fc8", x"7fc8", x"7fc8", x"7fc8", x"7fc8", 
    x"7fc7", x"7fc7", x"7fc7", x"7fc7", x"7fc7", x"7fc6", x"7fc6", x"7fc6", 
    x"7fc6", x"7fc6", x"7fc6", x"7fc5", x"7fc5", x"7fc5", x"7fc5", x"7fc5", 
    x"7fc4", x"7fc4", x"7fc4", x"7fc4", x"7fc4", x"7fc3", x"7fc3", x"7fc3", 
    x"7fc3", x"7fc3", x"7fc2", x"7fc2", x"7fc2", x"7fc2", x"7fc2", x"7fc2", 
    x"7fc1", x"7fc1", x"7fc1", x"7fc1", x"7fc1", x"7fc0", x"7fc0", x"7fc0", 
    x"7fc0", x"7fc0", x"7fbf", x"7fbf", x"7fbf", x"7fbf", x"7fbf", x"7fbe", 
    x"7fbe", x"7fbe", x"7fbe", x"7fbe", x"7fbd", x"7fbd", x"7fbd", x"7fbd", 
    x"7fbd", x"7fbc", x"7fbc", x"7fbc", x"7fbc", x"7fbc", x"7fbb", x"7fbb", 
    x"7fbb", x"7fbb", x"7fbb", x"7fba", x"7fba", x"7fba", x"7fba", x"7fba", 
    x"7fb9", x"7fb9", x"7fb9", x"7fb9", x"7fb9", x"7fb8", x"7fb8", x"7fb8", 
    x"7fb8", x"7fb8", x"7fb7", x"7fb7", x"7fb7", x"7fb7", x"7fb6", x"7fb6", 
    x"7fb6", x"7fb6", x"7fb6", x"7fb5", x"7fb5", x"7fb5", x"7fb5", x"7fb5", 
    x"7fb4", x"7fb4", x"7fb4", x"7fb4", x"7fb4", x"7fb3", x"7fb3", x"7fb3", 
    x"7fb3", x"7fb2", x"7fb2", x"7fb2", x"7fb2", x"7fb2", x"7fb1", x"7fb1", 
    x"7fb1", x"7fb1", x"7fb1", x"7fb0", x"7fb0", x"7fb0", x"7fb0", x"7faf", 
    x"7faf", x"7faf", x"7faf", x"7faf", x"7fae", x"7fae", x"7fae", x"7fae", 
    x"7fad", x"7fad", x"7fad", x"7fad", x"7fad", x"7fac", x"7fac", x"7fac", 
    x"7fac", x"7fab", x"7fab", x"7fab", x"7fab", x"7fab", x"7faa", x"7faa", 
    x"7faa", x"7faa", x"7fa9", x"7fa9", x"7fa9", x"7fa9", x"7fa9", x"7fa8", 
    x"7fa8", x"7fa8", x"7fa8", x"7fa7", x"7fa7", x"7fa7", x"7fa7", x"7fa6", 
    x"7fa6", x"7fa6", x"7fa6", x"7fa6", x"7fa5", x"7fa5", x"7fa5", x"7fa5", 
    x"7fa4", x"7fa4", x"7fa4", x"7fa4", x"7fa3", x"7fa3", x"7fa3", x"7fa3", 
    x"7fa2", x"7fa2", x"7fa2", x"7fa2", x"7fa2", x"7fa1", x"7fa1", x"7fa1", 
    x"7fa1", x"7fa0", x"7fa0", x"7fa0", x"7fa0", x"7f9f", x"7f9f", x"7f9f", 
    x"7f9f", x"7f9e", x"7f9e", x"7f9e", x"7f9e", x"7f9d", x"7f9d", x"7f9d", 
    x"7f9d", x"7f9c", x"7f9c", x"7f9c", x"7f9c", x"7f9c", x"7f9b", x"7f9b", 
    x"7f9b", x"7f9b", x"7f9a", x"7f9a", x"7f9a", x"7f9a", x"7f99", x"7f99", 
    x"7f99", x"7f99", x"7f98", x"7f98", x"7f98", x"7f98", x"7f97", x"7f97", 
    x"7f97", x"7f97", x"7f96", x"7f96", x"7f96", x"7f96", x"7f95", x"7f95", 
    x"7f95", x"7f95", x"7f94", x"7f94", x"7f94", x"7f94", x"7f93", x"7f93", 
    x"7f93", x"7f93", x"7f92", x"7f92", x"7f92", x"7f91", x"7f91", x"7f91", 
    x"7f91", x"7f90", x"7f90", x"7f90", x"7f90", x"7f8f", x"7f8f", x"7f8f", 
    x"7f8f", x"7f8e", x"7f8e", x"7f8e", x"7f8e", x"7f8d", x"7f8d", x"7f8d", 
    x"7f8d", x"7f8c", x"7f8c", x"7f8c", x"7f8c", x"7f8b", x"7f8b", x"7f8b", 
    x"7f8a", x"7f8a", x"7f8a", x"7f8a", x"7f89", x"7f89", x"7f89", x"7f89", 
    x"7f88", x"7f88", x"7f88", x"7f88", x"7f87", x"7f87", x"7f87", x"7f86", 
    x"7f86", x"7f86", x"7f86", x"7f85", x"7f85", x"7f85", x"7f85", x"7f84", 
    x"7f84", x"7f84", x"7f83", x"7f83", x"7f83", x"7f83", x"7f82", x"7f82", 
    x"7f82", x"7f82", x"7f81", x"7f81", x"7f81", x"7f80", x"7f80", x"7f80", 
    x"7f80", x"7f7f", x"7f7f", x"7f7f", x"7f7f", x"7f7e", x"7f7e", x"7f7e", 
    x"7f7d", x"7f7d", x"7f7d", x"7f7d", x"7f7c", x"7f7c", x"7f7c", x"7f7b", 
    x"7f7b", x"7f7b", x"7f7b", x"7f7a", x"7f7a", x"7f7a", x"7f79", x"7f79", 
    x"7f79", x"7f79", x"7f78", x"7f78", x"7f78", x"7f77", x"7f77", x"7f77", 
    x"7f77", x"7f76", x"7f76", x"7f76", x"7f75", x"7f75", x"7f75", x"7f75", 
    x"7f74", x"7f74", x"7f74", x"7f73", x"7f73", x"7f73", x"7f73", x"7f72", 
    x"7f72", x"7f72", x"7f71", x"7f71", x"7f71", x"7f71", x"7f70", x"7f70", 
    x"7f70", x"7f6f", x"7f6f", x"7f6f", x"7f6e", x"7f6e", x"7f6e", x"7f6e", 
    x"7f6d", x"7f6d", x"7f6d", x"7f6c", x"7f6c", x"7f6c", x"7f6c", x"7f6b", 
    x"7f6b", x"7f6b", x"7f6a", x"7f6a", x"7f6a", x"7f69", x"7f69", x"7f69", 
    x"7f69", x"7f68", x"7f68", x"7f68", x"7f67", x"7f67", x"7f67", x"7f66", 
    x"7f66", x"7f66", x"7f65", x"7f65", x"7f65", x"7f65", x"7f64", x"7f64", 
    x"7f64", x"7f63", x"7f63", x"7f63", x"7f62", x"7f62", x"7f62", x"7f62", 
    x"7f61", x"7f61", x"7f61", x"7f60", x"7f60", x"7f60", x"7f5f", x"7f5f", 
    x"7f5f", x"7f5e", x"7f5e", x"7f5e", x"7f5e", x"7f5d", x"7f5d", x"7f5d", 
    x"7f5c", x"7f5c", x"7f5c", x"7f5b", x"7f5b", x"7f5b", x"7f5a", x"7f5a", 
    x"7f5a", x"7f59", x"7f59", x"7f59", x"7f58", x"7f58", x"7f58", x"7f58", 
    x"7f57", x"7f57", x"7f57", x"7f56", x"7f56", x"7f56", x"7f55", x"7f55", 
    x"7f55", x"7f54", x"7f54", x"7f54", x"7f53", x"7f53", x"7f53", x"7f52", 
    x"7f52", x"7f52", x"7f51", x"7f51", x"7f51", x"7f50", x"7f50", x"7f50", 
    x"7f50", x"7f4f", x"7f4f", x"7f4f", x"7f4e", x"7f4e", x"7f4e", x"7f4d", 
    x"7f4d", x"7f4d", x"7f4c", x"7f4c", x"7f4c", x"7f4b", x"7f4b", x"7f4b", 
    x"7f4a", x"7f4a", x"7f4a", x"7f49", x"7f49", x"7f49", x"7f48", x"7f48", 
    x"7f48", x"7f47", x"7f47", x"7f47", x"7f46", x"7f46", x"7f46", x"7f45", 
    x"7f45", x"7f45", x"7f44", x"7f44", x"7f44", x"7f43", x"7f43", x"7f43", 
    x"7f42", x"7f42", x"7f42", x"7f41", x"7f41", x"7f41", x"7f40", x"7f40", 
    x"7f40", x"7f3f", x"7f3f", x"7f3f", x"7f3e", x"7f3e", x"7f3e", x"7f3d", 
    x"7f3d", x"7f3d", x"7f3c", x"7f3c", x"7f3b", x"7f3b", x"7f3b", x"7f3a", 
    x"7f3a", x"7f3a", x"7f39", x"7f39", x"7f39", x"7f38", x"7f38", x"7f38", 
    x"7f37", x"7f37", x"7f37", x"7f36", x"7f36", x"7f36", x"7f35", x"7f35", 
    x"7f35", x"7f34", x"7f34", x"7f34", x"7f33", x"7f33", x"7f32", x"7f32", 
    x"7f32", x"7f31", x"7f31", x"7f31", x"7f30", x"7f30", x"7f30", x"7f2f", 
    x"7f2f", x"7f2f", x"7f2e", x"7f2e", x"7f2e", x"7f2d", x"7f2d", x"7f2c", 
    x"7f2c", x"7f2c", x"7f2b", x"7f2b", x"7f2b", x"7f2a", x"7f2a", x"7f2a", 
    x"7f29", x"7f29", x"7f29", x"7f28", x"7f28", x"7f27", x"7f27", x"7f27", 
    x"7f26", x"7f26", x"7f26", x"7f25", x"7f25", x"7f25", x"7f24", x"7f24", 
    x"7f23", x"7f23", x"7f23", x"7f22", x"7f22", x"7f22", x"7f21", x"7f21", 
    x"7f21", x"7f20", x"7f20", x"7f1f", x"7f1f", x"7f1f", x"7f1e", x"7f1e", 
    x"7f1e", x"7f1d", x"7f1d", x"7f1d", x"7f1c", x"7f1c", x"7f1b", x"7f1b", 
    x"7f1b", x"7f1a", x"7f1a", x"7f1a", x"7f19", x"7f19", x"7f18", x"7f18", 
    x"7f18", x"7f17", x"7f17", x"7f17", x"7f16", x"7f16", x"7f15", x"7f15", 
    x"7f15", x"7f14", x"7f14", x"7f14", x"7f13", x"7f13", x"7f12", x"7f12", 
    x"7f12", x"7f11", x"7f11", x"7f11", x"7f10", x"7f10", x"7f0f", x"7f0f", 
    x"7f0f", x"7f0e", x"7f0e", x"7f0e", x"7f0d", x"7f0d", x"7f0c", x"7f0c", 
    x"7f0c", x"7f0b", x"7f0b", x"7f0a", x"7f0a", x"7f0a", x"7f09", x"7f09", 
    x"7f09", x"7f08", x"7f08", x"7f07", x"7f07", x"7f07", x"7f06", x"7f06", 
    x"7f05", x"7f05", x"7f05", x"7f04", x"7f04", x"7f04", x"7f03", x"7f03", 
    x"7f02", x"7f02", x"7f02", x"7f01", x"7f01", x"7f00", x"7f00", x"7f00", 
    x"7eff", x"7eff", x"7efe", x"7efe", x"7efe", x"7efd", x"7efd", x"7efd", 
    x"7efc", x"7efc", x"7efb", x"7efb", x"7efb", x"7efa", x"7efa", x"7ef9", 
    x"7ef9", x"7ef9", x"7ef8", x"7ef8", x"7ef7", x"7ef7", x"7ef7", x"7ef6", 
    x"7ef6", x"7ef5", x"7ef5", x"7ef5", x"7ef4", x"7ef4", x"7ef3", x"7ef3", 
    x"7ef3", x"7ef2", x"7ef2", x"7ef1", x"7ef1", x"7ef1", x"7ef0", x"7ef0", 
    x"7eef", x"7eef", x"7eef", x"7eee", x"7eee", x"7eed", x"7eed", x"7eed", 
    x"7eec", x"7eec", x"7eeb", x"7eeb", x"7eea", x"7eea", x"7eea", x"7ee9", 
    x"7ee9", x"7ee8", x"7ee8", x"7ee8", x"7ee7", x"7ee7", x"7ee6", x"7ee6", 
    x"7ee6", x"7ee5", x"7ee5", x"7ee4", x"7ee4", x"7ee4", x"7ee3", x"7ee3", 
    x"7ee2", x"7ee2", x"7ee1", x"7ee1", x"7ee1", x"7ee0", x"7ee0", x"7edf", 
    x"7edf", x"7edf", x"7ede", x"7ede", x"7edd", x"7edd", x"7edc", x"7edc", 
    x"7edc", x"7edb", x"7edb", x"7eda", x"7eda", x"7eda", x"7ed9", x"7ed9", 
    x"7ed8", x"7ed8", x"7ed7", x"7ed7", x"7ed7", x"7ed6", x"7ed6", x"7ed5", 
    x"7ed5", x"7ed4", x"7ed4", x"7ed4", x"7ed3", x"7ed3", x"7ed2", x"7ed2", 
    x"7ed2", x"7ed1", x"7ed1", x"7ed0", x"7ed0", x"7ecf", x"7ecf", x"7ecf", 
    x"7ece", x"7ece", x"7ecd", x"7ecd", x"7ecc", x"7ecc", x"7ecc", x"7ecb", 
    x"7ecb", x"7eca", x"7eca", x"7ec9", x"7ec9", x"7ec9", x"7ec8", x"7ec8", 
    x"7ec7", x"7ec7", x"7ec6", x"7ec6", x"7ec5", x"7ec5", x"7ec5", x"7ec4", 
    x"7ec4", x"7ec3", x"7ec3", x"7ec2", x"7ec2", x"7ec2", x"7ec1", x"7ec1", 
    x"7ec0", x"7ec0", x"7ebf", x"7ebf", x"7ebf", x"7ebe", x"7ebe", x"7ebd", 
    x"7ebd", x"7ebc", x"7ebc", x"7ebb", x"7ebb", x"7ebb", x"7eba", x"7eba", 
    x"7eb9", x"7eb9", x"7eb8", x"7eb8", x"7eb7", x"7eb7", x"7eb7", x"7eb6", 
    x"7eb6", x"7eb5", x"7eb5", x"7eb4", x"7eb4", x"7eb3", x"7eb3", x"7eb3", 
    x"7eb2", x"7eb2", x"7eb1", x"7eb1", x"7eb0", x"7eb0", x"7eaf", x"7eaf", 
    x"7eaf", x"7eae", x"7eae", x"7ead", x"7ead", x"7eac", x"7eac", x"7eab", 
    x"7eab", x"7eaa", x"7eaa", x"7eaa", x"7ea9", x"7ea9", x"7ea8", x"7ea8", 
    x"7ea7", x"7ea7", x"7ea6", x"7ea6", x"7ea6", x"7ea5", x"7ea5", x"7ea4", 
    x"7ea4", x"7ea3", x"7ea3", x"7ea2", x"7ea2", x"7ea1", x"7ea1", x"7ea0", 
    x"7ea0", x"7ea0", x"7e9f", x"7e9f", x"7e9e", x"7e9e", x"7e9d", x"7e9d", 
    x"7e9c", x"7e9c", x"7e9b", x"7e9b", x"7e9b", x"7e9a", x"7e9a", x"7e99", 
    x"7e99", x"7e98", x"7e98", x"7e97", x"7e97", x"7e96", x"7e96", x"7e95", 
    x"7e95", x"7e94", x"7e94", x"7e94", x"7e93", x"7e93", x"7e92", x"7e92", 
    x"7e91", x"7e91", x"7e90", x"7e90", x"7e8f", x"7e8f", x"7e8e", x"7e8e", 
    x"7e8d", x"7e8d", x"7e8d", x"7e8c", x"7e8c", x"7e8b", x"7e8b", x"7e8a", 
    x"7e8a", x"7e89", x"7e89", x"7e88", x"7e88", x"7e87", x"7e87", x"7e86", 
    x"7e86", x"7e85", x"7e85", x"7e84", x"7e84", x"7e83", x"7e83", x"7e83", 
    x"7e82", x"7e82", x"7e81", x"7e81", x"7e80", x"7e80", x"7e7f", x"7e7f", 
    x"7e7e", x"7e7e", x"7e7d", x"7e7d", x"7e7c", x"7e7c", x"7e7b", x"7e7b", 
    x"7e7a", x"7e7a", x"7e79", x"7e79", x"7e78", x"7e78", x"7e77", x"7e77", 
    x"7e77", x"7e76", x"7e76", x"7e75", x"7e75", x"7e74", x"7e74", x"7e73", 
    x"7e73", x"7e72", x"7e72", x"7e71", x"7e71", x"7e70", x"7e70", x"7e6f", 
    x"7e6f", x"7e6e", x"7e6e", x"7e6d", x"7e6d", x"7e6c", x"7e6c", x"7e6b", 
    x"7e6b", x"7e6a", x"7e6a", x"7e69", x"7e69", x"7e68", x"7e68", x"7e67", 
    x"7e67", x"7e66", x"7e66", x"7e65", x"7e65", x"7e64", x"7e64", x"7e63", 
    x"7e63", x"7e62", x"7e62", x"7e61", x"7e61", x"7e60", x"7e60", x"7e5f", 
    x"7e5f", x"7e5e", x"7e5e", x"7e5d", x"7e5d", x"7e5c", x"7e5c", x"7e5b", 
    x"7e5b", x"7e5a", x"7e5a", x"7e59", x"7e59", x"7e58", x"7e58", x"7e57", 
    x"7e57", x"7e56", x"7e56", x"7e55", x"7e55", x"7e54", x"7e54", x"7e53", 
    x"7e53", x"7e52", x"7e52", x"7e51", x"7e51", x"7e50", x"7e50", x"7e4f", 
    x"7e4f", x"7e4e", x"7e4e", x"7e4d", x"7e4d", x"7e4c", x"7e4c", x"7e4b", 
    x"7e4b", x"7e4a", x"7e4a", x"7e49", x"7e49", x"7e48", x"7e48", x"7e47", 
    x"7e47", x"7e46", x"7e46", x"7e45", x"7e45", x"7e44", x"7e44", x"7e43", 
    x"7e42", x"7e42", x"7e41", x"7e41", x"7e40", x"7e40", x"7e3f", x"7e3f", 
    x"7e3e", x"7e3e", x"7e3d", x"7e3d", x"7e3c", x"7e3c", x"7e3b", x"7e3b", 
    x"7e3a", x"7e3a", x"7e39", x"7e39", x"7e38", x"7e38", x"7e37", x"7e37", 
    x"7e36", x"7e36", x"7e35", x"7e34", x"7e34", x"7e33", x"7e33", x"7e32", 
    x"7e32", x"7e31", x"7e31", x"7e30", x"7e30", x"7e2f", x"7e2f", x"7e2e", 
    x"7e2e", x"7e2d", x"7e2d", x"7e2c", x"7e2c", x"7e2b", x"7e2a", x"7e2a", 
    x"7e29", x"7e29", x"7e28", x"7e28", x"7e27", x"7e27", x"7e26", x"7e26", 
    x"7e25", x"7e25", x"7e24", x"7e24", x"7e23", x"7e22", x"7e22", x"7e21", 
    x"7e21", x"7e20", x"7e20", x"7e1f", x"7e1f", x"7e1e", x"7e1e", x"7e1d", 
    x"7e1d", x"7e1c", x"7e1c", x"7e1b", x"7e1a", x"7e1a", x"7e19", x"7e19", 
    x"7e18", x"7e18", x"7e17", x"7e17", x"7e16", x"7e16", x"7e15", x"7e15", 
    x"7e14", x"7e13", x"7e13", x"7e12", x"7e12", x"7e11", x"7e11", x"7e10", 
    x"7e10", x"7e0f", x"7e0f", x"7e0e", x"7e0d", x"7e0d", x"7e0c", x"7e0c", 
    x"7e0b", x"7e0b", x"7e0a", x"7e0a", x"7e09", x"7e09", x"7e08", x"7e07", 
    x"7e07", x"7e06", x"7e06", x"7e05", x"7e05", x"7e04", x"7e04", x"7e03", 
    x"7e02", x"7e02", x"7e01", x"7e01", x"7e00", x"7e00", x"7dff", x"7dff", 
    x"7dfe", x"7dfd", x"7dfd", x"7dfc", x"7dfc", x"7dfb", x"7dfb", x"7dfa", 
    x"7dfa", x"7df9", x"7df8", x"7df8", x"7df7", x"7df7", x"7df6", x"7df6", 
    x"7df5", x"7df5", x"7df4", x"7df3", x"7df3", x"7df2", x"7df2", x"7df1", 
    x"7df1", x"7df0", x"7df0", x"7def", x"7dee", x"7dee", x"7ded", x"7ded", 
    x"7dec", x"7dec", x"7deb", x"7dea", x"7dea", x"7de9", x"7de9", x"7de8", 
    x"7de8", x"7de7", x"7de7", x"7de6", x"7de5", x"7de5", x"7de4", x"7de4", 
    x"7de3", x"7de3", x"7de2", x"7de1", x"7de1", x"7de0", x"7de0", x"7ddf", 
    x"7ddf", x"7dde", x"7ddd", x"7ddd", x"7ddc", x"7ddc", x"7ddb", x"7ddb", 
    x"7dda", x"7dd9", x"7dd9", x"7dd8", x"7dd8", x"7dd7", x"7dd7", x"7dd6", 
    x"7dd5", x"7dd5", x"7dd4", x"7dd4", x"7dd3", x"7dd3", x"7dd2", x"7dd1", 
    x"7dd1", x"7dd0", x"7dd0", x"7dcf", x"7dce", x"7dce", x"7dcd", x"7dcd", 
    x"7dcc", x"7dcc", x"7dcb", x"7dca", x"7dca", x"7dc9", x"7dc9", x"7dc8", 
    x"7dc8", x"7dc7", x"7dc6", x"7dc6", x"7dc5", x"7dc5", x"7dc4", x"7dc3", 
    x"7dc3", x"7dc2", x"7dc2", x"7dc1", x"7dc1", x"7dc0", x"7dbf", x"7dbf", 
    x"7dbe", x"7dbe", x"7dbd", x"7dbc", x"7dbc", x"7dbb", x"7dbb", x"7dba", 
    x"7db9", x"7db9", x"7db8", x"7db8", x"7db7", x"7db7", x"7db6", x"7db5", 
    x"7db5", x"7db4", x"7db4", x"7db3", x"7db2", x"7db2", x"7db1", x"7db1", 
    x"7db0", x"7daf", x"7daf", x"7dae", x"7dae", x"7dad", x"7dac", x"7dac", 
    x"7dab", x"7dab", x"7daa", x"7da9", x"7da9", x"7da8", x"7da8", x"7da7", 
    x"7da6", x"7da6", x"7da5", x"7da5", x"7da4", x"7da3", x"7da3", x"7da2", 
    x"7da2", x"7da1", x"7da0", x"7da0", x"7d9f", x"7d9f", x"7d9e", x"7d9d", 
    x"7d9d", x"7d9c", x"7d9c", x"7d9b", x"7d9a", x"7d9a", x"7d99", x"7d99", 
    x"7d98", x"7d97", x"7d97", x"7d96", x"7d96", x"7d95", x"7d94", x"7d94", 
    x"7d93", x"7d93", x"7d92", x"7d91", x"7d91", x"7d90", x"7d90", x"7d8f", 
    x"7d8e", x"7d8e", x"7d8d", x"7d8c", x"7d8c", x"7d8b", x"7d8b", x"7d8a", 
    x"7d89", x"7d89", x"7d88", x"7d88", x"7d87", x"7d86", x"7d86", x"7d85", 
    x"7d84", x"7d84", x"7d83", x"7d83", x"7d82", x"7d81", x"7d81", x"7d80", 
    x"7d80", x"7d7f", x"7d7e", x"7d7e", x"7d7d", x"7d7c", x"7d7c", x"7d7b", 
    x"7d7b", x"7d7a", x"7d79", x"7d79", x"7d78", x"7d77", x"7d77", x"7d76", 
    x"7d76", x"7d75", x"7d74", x"7d74", x"7d73", x"7d73", x"7d72", x"7d71", 
    x"7d71", x"7d70", x"7d6f", x"7d6f", x"7d6e", x"7d6e", x"7d6d", x"7d6c", 
    x"7d6c", x"7d6b", x"7d6a", x"7d6a", x"7d69", x"7d68", x"7d68", x"7d67", 
    x"7d67", x"7d66", x"7d65", x"7d65", x"7d64", x"7d63", x"7d63", x"7d62", 
    x"7d62", x"7d61", x"7d60", x"7d60", x"7d5f", x"7d5e", x"7d5e", x"7d5d", 
    x"7d5c", x"7d5c", x"7d5b", x"7d5b", x"7d5a", x"7d59", x"7d59", x"7d58", 
    x"7d57", x"7d57", x"7d56", x"7d56", x"7d55", x"7d54", x"7d54", x"7d53", 
    x"7d52", x"7d52", x"7d51", x"7d50", x"7d50", x"7d4f", x"7d4e", x"7d4e", 
    x"7d4d", x"7d4d", x"7d4c", x"7d4b", x"7d4b", x"7d4a", x"7d49", x"7d49", 
    x"7d48", x"7d47", x"7d47", x"7d46", x"7d45", x"7d45", x"7d44", x"7d44", 
    x"7d43", x"7d42", x"7d42", x"7d41", x"7d40", x"7d40", x"7d3f", x"7d3e", 
    x"7d3e", x"7d3d", x"7d3c", x"7d3c", x"7d3b", x"7d3a", x"7d3a", x"7d39", 
    x"7d39", x"7d38", x"7d37", x"7d37", x"7d36", x"7d35", x"7d35", x"7d34", 
    x"7d33", x"7d33", x"7d32", x"7d31", x"7d31", x"7d30", x"7d2f", x"7d2f", 
    x"7d2e", x"7d2d", x"7d2d", x"7d2c", x"7d2b", x"7d2b", x"7d2a", x"7d29", 
    x"7d29", x"7d28", x"7d28", x"7d27", x"7d26", x"7d26", x"7d25", x"7d24", 
    x"7d24", x"7d23", x"7d22", x"7d22", x"7d21", x"7d20", x"7d20", x"7d1f", 
    x"7d1e", x"7d1e", x"7d1d", x"7d1c", x"7d1c", x"7d1b", x"7d1a", x"7d1a", 
    x"7d19", x"7d18", x"7d18", x"7d17", x"7d16", x"7d16", x"7d15", x"7d14", 
    x"7d14", x"7d13", x"7d12", x"7d12", x"7d11", x"7d10", x"7d10", x"7d0f", 
    x"7d0e", x"7d0e", x"7d0d", x"7d0c", x"7d0c", x"7d0b", x"7d0a", x"7d0a", 
    x"7d09", x"7d08", x"7d08", x"7d07", x"7d06", x"7d06", x"7d05", x"7d04", 
    x"7d04", x"7d03", x"7d02", x"7d02", x"7d01", x"7d00", x"7cff", x"7cff", 
    x"7cfe", x"7cfd", x"7cfd", x"7cfc", x"7cfb", x"7cfb", x"7cfa", x"7cf9", 
    x"7cf9", x"7cf8", x"7cf7", x"7cf7", x"7cf6", x"7cf5", x"7cf5", x"7cf4", 
    x"7cf3", x"7cf3", x"7cf2", x"7cf1", x"7cf1", x"7cf0", x"7cef", x"7cee", 
    x"7cee", x"7ced", x"7cec", x"7cec", x"7ceb", x"7cea", x"7cea", x"7ce9", 
    x"7ce8", x"7ce8", x"7ce7", x"7ce6", x"7ce6", x"7ce5", x"7ce4", x"7ce4", 
    x"7ce3", x"7ce2", x"7ce1", x"7ce1", x"7ce0", x"7cdf", x"7cdf", x"7cde", 
    x"7cdd", x"7cdd", x"7cdc", x"7cdb", x"7cdb", x"7cda", x"7cd9", x"7cd8", 
    x"7cd8", x"7cd7", x"7cd6", x"7cd6", x"7cd5", x"7cd4", x"7cd4", x"7cd3", 
    x"7cd2", x"7cd2", x"7cd1", x"7cd0", x"7ccf", x"7ccf", x"7cce", x"7ccd", 
    x"7ccd", x"7ccc", x"7ccb", x"7ccb", x"7cca", x"7cc9", x"7cc8", x"7cc8", 
    x"7cc7", x"7cc6", x"7cc6", x"7cc5", x"7cc4", x"7cc4", x"7cc3", x"7cc2", 
    x"7cc1", x"7cc1", x"7cc0", x"7cbf", x"7cbf", x"7cbe", x"7cbd", x"7cbd", 
    x"7cbc", x"7cbb", x"7cba", x"7cba", x"7cb9", x"7cb8", x"7cb8", x"7cb7", 
    x"7cb6", x"7cb5", x"7cb5", x"7cb4", x"7cb3", x"7cb3", x"7cb2", x"7cb1", 
    x"7cb1", x"7cb0", x"7caf", x"7cae", x"7cae", x"7cad", x"7cac", x"7cac", 
    x"7cab", x"7caa", x"7ca9", x"7ca9", x"7ca8", x"7ca7", x"7ca7", x"7ca6", 
    x"7ca5", x"7ca4", x"7ca4", x"7ca3", x"7ca2", x"7ca2", x"7ca1", x"7ca0", 
    x"7c9f", x"7c9f", x"7c9e", x"7c9d", x"7c9d", x"7c9c", x"7c9b", x"7c9a", 
    x"7c9a", x"7c99", x"7c98", x"7c98", x"7c97", x"7c96", x"7c95", x"7c95", 
    x"7c94", x"7c93", x"7c92", x"7c92", x"7c91", x"7c90", x"7c90", x"7c8f", 
    x"7c8e", x"7c8d", x"7c8d", x"7c8c", x"7c8b", x"7c8a", x"7c8a", x"7c89", 
    x"7c88", x"7c88", x"7c87", x"7c86", x"7c85", x"7c85", x"7c84", x"7c83", 
    x"7c83", x"7c82", x"7c81", x"7c80", x"7c80", x"7c7f", x"7c7e", x"7c7d", 
    x"7c7d", x"7c7c", x"7c7b", x"7c7a", x"7c7a", x"7c79", x"7c78", x"7c78", 
    x"7c77", x"7c76", x"7c75", x"7c75", x"7c74", x"7c73", x"7c72", x"7c72", 
    x"7c71", x"7c70", x"7c6f", x"7c6f", x"7c6e", x"7c6d", x"7c6d", x"7c6c", 
    x"7c6b", x"7c6a", x"7c6a", x"7c69", x"7c68", x"7c67", x"7c67", x"7c66", 
    x"7c65", x"7c64", x"7c64", x"7c63", x"7c62", x"7c61", x"7c61", x"7c60", 
    x"7c5f", x"7c5e", x"7c5e", x"7c5d", x"7c5c", x"7c5c", x"7c5b", x"7c5a", 
    x"7c59", x"7c59", x"7c58", x"7c57", x"7c56", x"7c56", x"7c55", x"7c54", 
    x"7c53", x"7c53", x"7c52", x"7c51", x"7c50", x"7c50", x"7c4f", x"7c4e", 
    x"7c4d", x"7c4d", x"7c4c", x"7c4b", x"7c4a", x"7c4a", x"7c49", x"7c48", 
    x"7c47", x"7c47", x"7c46", x"7c45", x"7c44", x"7c44", x"7c43", x"7c42", 
    x"7c41", x"7c41", x"7c40", x"7c3f", x"7c3e", x"7c3e", x"7c3d", x"7c3c", 
    x"7c3b", x"7c3a", x"7c3a", x"7c39", x"7c38", x"7c37", x"7c37", x"7c36", 
    x"7c35", x"7c34", x"7c34", x"7c33", x"7c32", x"7c31", x"7c31", x"7c30", 
    x"7c2f", x"7c2e", x"7c2e", x"7c2d", x"7c2c", x"7c2b", x"7c2b", x"7c2a", 
    x"7c29", x"7c28", x"7c27", x"7c27", x"7c26", x"7c25", x"7c24", x"7c24", 
    x"7c23", x"7c22", x"7c21", x"7c21", x"7c20", x"7c1f", x"7c1e", x"7c1e", 
    x"7c1d", x"7c1c", x"7c1b", x"7c1a", x"7c1a", x"7c19", x"7c18", x"7c17", 
    x"7c17", x"7c16", x"7c15", x"7c14", x"7c14", x"7c13", x"7c12", x"7c11", 
    x"7c10", x"7c10", x"7c0f", x"7c0e", x"7c0d", x"7c0d", x"7c0c", x"7c0b", 
    x"7c0a", x"7c09", x"7c09", x"7c08", x"7c07", x"7c06", x"7c06", x"7c05", 
    x"7c04", x"7c03", x"7c02", x"7c02", x"7c01", x"7c00", x"7bff", x"7bff", 
    x"7bfe", x"7bfd", x"7bfc", x"7bfb", x"7bfb", x"7bfa", x"7bf9", x"7bf8", 
    x"7bf8", x"7bf7", x"7bf6", x"7bf5", x"7bf4", x"7bf4", x"7bf3", x"7bf2", 
    x"7bf1", x"7bf1", x"7bf0", x"7bef", x"7bee", x"7bed", x"7bed", x"7bec", 
    x"7beb", x"7bea", x"7be9", x"7be9", x"7be8", x"7be7", x"7be6", x"7be6", 
    x"7be5", x"7be4", x"7be3", x"7be2", x"7be2", x"7be1", x"7be0", x"7bdf", 
    x"7bde", x"7bde", x"7bdd", x"7bdc", x"7bdb", x"7bda", x"7bda", x"7bd9", 
    x"7bd8", x"7bd7", x"7bd6", x"7bd6", x"7bd5", x"7bd4", x"7bd3", x"7bd2", 
    x"7bd2", x"7bd1", x"7bd0", x"7bcf", x"7bcf", x"7bce", x"7bcd", x"7bcc", 
    x"7bcb", x"7bcb", x"7bca", x"7bc9", x"7bc8", x"7bc7", x"7bc7", x"7bc6", 
    x"7bc5", x"7bc4", x"7bc3", x"7bc3", x"7bc2", x"7bc1", x"7bc0", x"7bbf", 
    x"7bbf", x"7bbe", x"7bbd", x"7bbc", x"7bbb", x"7bba", x"7bba", x"7bb9", 
    x"7bb8", x"7bb7", x"7bb6", x"7bb6", x"7bb5", x"7bb4", x"7bb3", x"7bb2", 
    x"7bb2", x"7bb1", x"7bb0", x"7baf", x"7bae", x"7bae", x"7bad", x"7bac", 
    x"7bab", x"7baa", x"7baa", x"7ba9", x"7ba8", x"7ba7", x"7ba6", x"7ba5", 
    x"7ba5", x"7ba4", x"7ba3", x"7ba2", x"7ba1", x"7ba1", x"7ba0", x"7b9f", 
    x"7b9e", x"7b9d", x"7b9d", x"7b9c", x"7b9b", x"7b9a", x"7b99", x"7b98", 
    x"7b98", x"7b97", x"7b96", x"7b95", x"7b94", x"7b94", x"7b93", x"7b92", 
    x"7b91", x"7b90", x"7b8f", x"7b8f", x"7b8e", x"7b8d", x"7b8c", x"7b8b", 
    x"7b8b", x"7b8a", x"7b89", x"7b88", x"7b87", x"7b86", x"7b86", x"7b85", 
    x"7b84", x"7b83", x"7b82", x"7b81", x"7b81", x"7b80", x"7b7f", x"7b7e", 
    x"7b7d", x"7b7d", x"7b7c", x"7b7b", x"7b7a", x"7b79", x"7b78", x"7b78", 
    x"7b77", x"7b76", x"7b75", x"7b74", x"7b73", x"7b73", x"7b72", x"7b71", 
    x"7b70", x"7b6f", x"7b6e", x"7b6e", x"7b6d", x"7b6c", x"7b6b", x"7b6a", 
    x"7b69", x"7b69", x"7b68", x"7b67", x"7b66", x"7b65", x"7b64", x"7b64", 
    x"7b63", x"7b62", x"7b61", x"7b60", x"7b5f", x"7b5f", x"7b5e", x"7b5d", 
    x"7b5c", x"7b5b", x"7b5a", x"7b5a", x"7b59", x"7b58", x"7b57", x"7b56", 
    x"7b55", x"7b54", x"7b54", x"7b53", x"7b52", x"7b51", x"7b50", x"7b4f", 
    x"7b4f", x"7b4e", x"7b4d", x"7b4c", x"7b4b", x"7b4a", x"7b4a", x"7b49", 
    x"7b48", x"7b47", x"7b46", x"7b45", x"7b44", x"7b44", x"7b43", x"7b42", 
    x"7b41", x"7b40", x"7b3f", x"7b3f", x"7b3e", x"7b3d", x"7b3c", x"7b3b", 
    x"7b3a", x"7b39", x"7b39", x"7b38", x"7b37", x"7b36", x"7b35", x"7b34", 
    x"7b33", x"7b33", x"7b32", x"7b31", x"7b30", x"7b2f", x"7b2e", x"7b2e", 
    x"7b2d", x"7b2c", x"7b2b", x"7b2a", x"7b29", x"7b28", x"7b28", x"7b27", 
    x"7b26", x"7b25", x"7b24", x"7b23", x"7b22", x"7b22", x"7b21", x"7b20", 
    x"7b1f", x"7b1e", x"7b1d", x"7b1c", x"7b1c", x"7b1b", x"7b1a", x"7b19", 
    x"7b18", x"7b17", x"7b16", x"7b16", x"7b15", x"7b14", x"7b13", x"7b12", 
    x"7b11", x"7b10", x"7b0f", x"7b0f", x"7b0e", x"7b0d", x"7b0c", x"7b0b", 
    x"7b0a", x"7b09", x"7b09", x"7b08", x"7b07", x"7b06", x"7b05", x"7b04", 
    x"7b03", x"7b02", x"7b02", x"7b01", x"7b00", x"7aff", x"7afe", x"7afd", 
    x"7afc", x"7afc", x"7afb", x"7afa", x"7af9", x"7af8", x"7af7", x"7af6", 
    x"7af5", x"7af5", x"7af4", x"7af3", x"7af2", x"7af1", x"7af0", x"7aef", 
    x"7aee", x"7aee", x"7aed", x"7aec", x"7aeb", x"7aea", x"7ae9", x"7ae8", 
    x"7ae7", x"7ae7", x"7ae6", x"7ae5", x"7ae4", x"7ae3", x"7ae2", x"7ae1", 
    x"7ae0", x"7ae0", x"7adf", x"7ade", x"7add", x"7adc", x"7adb", x"7ada", 
    x"7ad9", x"7ad8", x"7ad8", x"7ad7", x"7ad6", x"7ad5", x"7ad4", x"7ad3", 
    x"7ad2", x"7ad1", x"7ad1", x"7ad0", x"7acf", x"7ace", x"7acd", x"7acc", 
    x"7acb", x"7aca", x"7ac9", x"7ac9", x"7ac8", x"7ac7", x"7ac6", x"7ac5", 
    x"7ac4", x"7ac3", x"7ac2", x"7ac1", x"7ac1", x"7ac0", x"7abf", x"7abe", 
    x"7abd", x"7abc", x"7abb", x"7aba", x"7ab9", x"7ab9", x"7ab8", x"7ab7", 
    x"7ab6", x"7ab5", x"7ab4", x"7ab3", x"7ab2", x"7ab1", x"7ab0", x"7ab0", 
    x"7aaf", x"7aae", x"7aad", x"7aac", x"7aab", x"7aaa", x"7aa9", x"7aa8", 
    x"7aa8", x"7aa7", x"7aa6", x"7aa5", x"7aa4", x"7aa3", x"7aa2", x"7aa1", 
    x"7aa0", x"7a9f", x"7a9f", x"7a9e", x"7a9d", x"7a9c", x"7a9b", x"7a9a", 
    x"7a99", x"7a98", x"7a97", x"7a96", x"7a95", x"7a95", x"7a94", x"7a93", 
    x"7a92", x"7a91", x"7a90", x"7a8f", x"7a8e", x"7a8d", x"7a8c", x"7a8c", 
    x"7a8b", x"7a8a", x"7a89", x"7a88", x"7a87", x"7a86", x"7a85", x"7a84", 
    x"7a83", x"7a82", x"7a82", x"7a81", x"7a80", x"7a7f", x"7a7e", x"7a7d", 
    x"7a7c", x"7a7b", x"7a7a", x"7a79", x"7a78", x"7a78", x"7a77", x"7a76", 
    x"7a75", x"7a74", x"7a73", x"7a72", x"7a71", x"7a70", x"7a6f", x"7a6e", 
    x"7a6d", x"7a6d", x"7a6c", x"7a6b", x"7a6a", x"7a69", x"7a68", x"7a67", 
    x"7a66", x"7a65", x"7a64", x"7a63", x"7a62", x"7a61", x"7a61", x"7a60", 
    x"7a5f", x"7a5e", x"7a5d", x"7a5c", x"7a5b", x"7a5a", x"7a59", x"7a58", 
    x"7a57", x"7a56", x"7a56", x"7a55", x"7a54", x"7a53", x"7a52", x"7a51", 
    x"7a50", x"7a4f", x"7a4e", x"7a4d", x"7a4c", x"7a4b", x"7a4a", x"7a49", 
    x"7a49", x"7a48", x"7a47", x"7a46", x"7a45", x"7a44", x"7a43", x"7a42", 
    x"7a41", x"7a40", x"7a3f", x"7a3e", x"7a3d", x"7a3c", x"7a3c", x"7a3b", 
    x"7a3a", x"7a39", x"7a38", x"7a37", x"7a36", x"7a35", x"7a34", x"7a33", 
    x"7a32", x"7a31", x"7a30", x"7a2f", x"7a2e", x"7a2e", x"7a2d", x"7a2c", 
    x"7a2b", x"7a2a", x"7a29", x"7a28", x"7a27", x"7a26", x"7a25", x"7a24", 
    x"7a23", x"7a22", x"7a21", x"7a20", x"7a1f", x"7a1e", x"7a1e", x"7a1d", 
    x"7a1c", x"7a1b", x"7a1a", x"7a19", x"7a18", x"7a17", x"7a16", x"7a15", 
    x"7a14", x"7a13", x"7a12", x"7a11", x"7a10", x"7a0f", x"7a0e", x"7a0e", 
    x"7a0d", x"7a0c", x"7a0b", x"7a0a", x"7a09", x"7a08", x"7a07", x"7a06", 
    x"7a05", x"7a04", x"7a03", x"7a02", x"7a01", x"7a00", x"79ff", x"79fe", 
    x"79fd", x"79fc", x"79fb", x"79fb", x"79fa", x"79f9", x"79f8", x"79f7", 
    x"79f6", x"79f5", x"79f4", x"79f3", x"79f2", x"79f1", x"79f0", x"79ef", 
    x"79ee", x"79ed", x"79ec", x"79eb", x"79ea", x"79e9", x"79e8", x"79e7", 
    x"79e6", x"79e6", x"79e5", x"79e4", x"79e3", x"79e2", x"79e1", x"79e0", 
    x"79df", x"79de", x"79dd", x"79dc", x"79db", x"79da", x"79d9", x"79d8", 
    x"79d7", x"79d6", x"79d5", x"79d4", x"79d3", x"79d2", x"79d1", x"79d0", 
    x"79cf", x"79ce", x"79cd", x"79cd", x"79cc", x"79cb", x"79ca", x"79c9", 
    x"79c8", x"79c7", x"79c6", x"79c5", x"79c4", x"79c3", x"79c2", x"79c1", 
    x"79c0", x"79bf", x"79be", x"79bd", x"79bc", x"79bb", x"79ba", x"79b9", 
    x"79b8", x"79b7", x"79b6", x"79b5", x"79b4", x"79b3", x"79b2", x"79b1", 
    x"79b0", x"79af", x"79ae", x"79ad", x"79ac", x"79ac", x"79ab", x"79aa", 
    x"79a9", x"79a8", x"79a7", x"79a6", x"79a5", x"79a4", x"79a3", x"79a2", 
    x"79a1", x"79a0", x"799f", x"799e", x"799d", x"799c", x"799b", x"799a", 
    x"7999", x"7998", x"7997", x"7996", x"7995", x"7994", x"7993", x"7992", 
    x"7991", x"7990", x"798f", x"798e", x"798d", x"798c", x"798b", x"798a", 
    x"7989", x"7988", x"7987", x"7986", x"7985", x"7984", x"7983", x"7982", 
    x"7981", x"7980", x"797f", x"797e", x"797d", x"797c", x"797b", x"797a", 
    x"7979", x"7978", x"7977", x"7976", x"7975", x"7974", x"7973", x"7972", 
    x"7971", x"7970", x"796f", x"796e", x"796d", x"796c", x"796b", x"796b", 
    x"796a", x"7969", x"7968", x"7967", x"7966", x"7965", x"7964", x"7963", 
    x"7962", x"7961", x"7960", x"795f", x"795e", x"795d", x"795c", x"795b", 
    x"795a", x"7959", x"7958", x"7957", x"7956", x"7955", x"7954", x"7953", 
    x"7952", x"7951", x"7950", x"794f", x"794e", x"794d", x"794c", x"794b", 
    x"794a", x"7949", x"7948", x"7947", x"7946", x"7945", x"7944", x"7943", 
    x"7941", x"7940", x"793f", x"793e", x"793d", x"793c", x"793b", x"793a", 
    x"7939", x"7938", x"7937", x"7936", x"7935", x"7934", x"7933", x"7932", 
    x"7931", x"7930", x"792f", x"792e", x"792d", x"792c", x"792b", x"792a", 
    x"7929", x"7928", x"7927", x"7926", x"7925", x"7924", x"7923", x"7922", 
    x"7921", x"7920", x"791f", x"791e", x"791d", x"791c", x"791b", x"791a", 
    x"7919", x"7918", x"7917", x"7916", x"7915", x"7914", x"7913", x"7912", 
    x"7911", x"7910", x"790f", x"790e", x"790d", x"790c", x"790b", x"790a", 
    x"7909", x"7908", x"7907", x"7906", x"7905", x"7904", x"7903", x"7902", 
    x"7901", x"7900", x"78fe", x"78fd", x"78fc", x"78fb", x"78fa", x"78f9", 
    x"78f8", x"78f7", x"78f6", x"78f5", x"78f4", x"78f3", x"78f2", x"78f1", 
    x"78f0", x"78ef", x"78ee", x"78ed", x"78ec", x"78eb", x"78ea", x"78e9", 
    x"78e8", x"78e7", x"78e6", x"78e5", x"78e4", x"78e3", x"78e2", x"78e1", 
    x"78e0", x"78df", x"78de", x"78dd", x"78db", x"78da", x"78d9", x"78d8", 
    x"78d7", x"78d6", x"78d5", x"78d4", x"78d3", x"78d2", x"78d1", x"78d0", 
    x"78cf", x"78ce", x"78cd", x"78cc", x"78cb", x"78ca", x"78c9", x"78c8", 
    x"78c7", x"78c6", x"78c5", x"78c4", x"78c3", x"78c2", x"78c0", x"78bf", 
    x"78be", x"78bd", x"78bc", x"78bb", x"78ba", x"78b9", x"78b8", x"78b7", 
    x"78b6", x"78b5", x"78b4", x"78b3", x"78b2", x"78b1", x"78b0", x"78af", 
    x"78ae", x"78ad", x"78ac", x"78ab", x"78a9", x"78a8", x"78a7", x"78a6", 
    x"78a5", x"78a4", x"78a3", x"78a2", x"78a1", x"78a0", x"789f", x"789e", 
    x"789d", x"789c", x"789b", x"789a", x"7899", x"7898", x"7897", x"7896", 
    x"7894", x"7893", x"7892", x"7891", x"7890", x"788f", x"788e", x"788d", 
    x"788c", x"788b", x"788a", x"7889", x"7888", x"7887", x"7886", x"7885", 
    x"7884", x"7883", x"7881", x"7880", x"787f", x"787e", x"787d", x"787c", 
    x"787b", x"787a", x"7879", x"7878", x"7877", x"7876", x"7875", x"7874", 
    x"7873", x"7872", x"7870", x"786f", x"786e", x"786d", x"786c", x"786b", 
    x"786a", x"7869", x"7868", x"7867", x"7866", x"7865", x"7864", x"7863", 
    x"7862", x"7860", x"785f", x"785e", x"785d", x"785c", x"785b", x"785a", 
    x"7859", x"7858", x"7857", x"7856", x"7855", x"7854", x"7853", x"7852", 
    x"7850", x"784f", x"784e", x"784d", x"784c", x"784b", x"784a", x"7849", 
    x"7848", x"7847", x"7846", x"7845", x"7844", x"7842", x"7841", x"7840", 
    x"783f", x"783e", x"783d", x"783c", x"783b", x"783a", x"7839", x"7838", 
    x"7837", x"7836", x"7834", x"7833", x"7832", x"7831", x"7830", x"782f", 
    x"782e", x"782d", x"782c", x"782b", x"782a", x"7829", x"7828", x"7826", 
    x"7825", x"7824", x"7823", x"7822", x"7821", x"7820", x"781f", x"781e", 
    x"781d", x"781c", x"781a", x"7819", x"7818", x"7817", x"7816", x"7815", 
    x"7814", x"7813", x"7812", x"7811", x"7810", x"780f", x"780d", x"780c", 
    x"780b", x"780a", x"7809", x"7808", x"7807", x"7806", x"7805", x"7804", 
    x"7803", x"7801", x"7800", x"77ff", x"77fe", x"77fd", x"77fc", x"77fb", 
    x"77fa", x"77f9", x"77f8", x"77f7", x"77f5", x"77f4", x"77f3", x"77f2", 
    x"77f1", x"77f0", x"77ef", x"77ee", x"77ed", x"77ec", x"77ea", x"77e9", 
    x"77e8", x"77e7", x"77e6", x"77e5", x"77e4", x"77e3", x"77e2", x"77e1", 
    x"77df", x"77de", x"77dd", x"77dc", x"77db", x"77da", x"77d9", x"77d8", 
    x"77d7", x"77d6", x"77d4", x"77d3", x"77d2", x"77d1", x"77d0", x"77cf", 
    x"77ce", x"77cd", x"77cc", x"77ca", x"77c9", x"77c8", x"77c7", x"77c6", 
    x"77c5", x"77c4", x"77c3", x"77c2", x"77c0", x"77bf", x"77be", x"77bd", 
    x"77bc", x"77bb", x"77ba", x"77b9", x"77b8", x"77b6", x"77b5", x"77b4", 
    x"77b3", x"77b2", x"77b1", x"77b0", x"77af", x"77ae", x"77ac", x"77ab", 
    x"77aa", x"77a9", x"77a8", x"77a7", x"77a6", x"77a5", x"77a4", x"77a2", 
    x"77a1", x"77a0", x"779f", x"779e", x"779d", x"779c", x"779b", x"7799", 
    x"7798", x"7797", x"7796", x"7795", x"7794", x"7793", x"7792", x"7791", 
    x"778f", x"778e", x"778d", x"778c", x"778b", x"778a", x"7789", x"7788", 
    x"7786", x"7785", x"7784", x"7783", x"7782", x"7781", x"7780", x"777f", 
    x"777d", x"777c", x"777b", x"777a", x"7779", x"7778", x"7777", x"7776", 
    x"7774", x"7773", x"7772", x"7771", x"7770", x"776f", x"776e", x"776d", 
    x"776b", x"776a", x"7769", x"7768", x"7767", x"7766", x"7765", x"7763", 
    x"7762", x"7761", x"7760", x"775f", x"775e", x"775d", x"775c", x"775a", 
    x"7759", x"7758", x"7757", x"7756", x"7755", x"7754", x"7752", x"7751", 
    x"7750", x"774f", x"774e", x"774d", x"774c", x"774a", x"7749", x"7748", 
    x"7747", x"7746", x"7745", x"7744", x"7742", x"7741", x"7740", x"773f", 
    x"773e", x"773d", x"773c", x"773a", x"7739", x"7738", x"7737", x"7736", 
    x"7735", x"7734", x"7732", x"7731", x"7730", x"772f", x"772e", x"772d", 
    x"772c", x"772a", x"7729", x"7728", x"7727", x"7726", x"7725", x"7724", 
    x"7722", x"7721", x"7720", x"771f", x"771e", x"771d", x"771c", x"771a", 
    x"7719", x"7718", x"7717", x"7716", x"7715", x"7713", x"7712", x"7711", 
    x"7710", x"770f", x"770e", x"770d", x"770b", x"770a", x"7709", x"7708", 
    x"7707", x"7706", x"7704", x"7703", x"7702", x"7701", x"7700", x"76ff", 
    x"76fe", x"76fc", x"76fb", x"76fa", x"76f9", x"76f8", x"76f7", x"76f5", 
    x"76f4", x"76f3", x"76f2", x"76f1", x"76f0", x"76ee", x"76ed", x"76ec", 
    x"76eb", x"76ea", x"76e9", x"76e7", x"76e6", x"76e5", x"76e4", x"76e3", 
    x"76e2", x"76e1", x"76df", x"76de", x"76dd", x"76dc", x"76db", x"76da", 
    x"76d8", x"76d7", x"76d6", x"76d5", x"76d4", x"76d3", x"76d1", x"76d0", 
    x"76cf", x"76ce", x"76cd", x"76cc", x"76ca", x"76c9", x"76c8", x"76c7", 
    x"76c6", x"76c4", x"76c3", x"76c2", x"76c1", x"76c0", x"76bf", x"76bd", 
    x"76bc", x"76bb", x"76ba", x"76b9", x"76b8", x"76b6", x"76b5", x"76b4", 
    x"76b3", x"76b2", x"76b1", x"76af", x"76ae", x"76ad", x"76ac", x"76ab", 
    x"76a9", x"76a8", x"76a7", x"76a6", x"76a5", x"76a4", x"76a2", x"76a1", 
    x"76a0", x"769f", x"769e", x"769d", x"769b", x"769a", x"7699", x"7698", 
    x"7697", x"7695", x"7694", x"7693", x"7692", x"7691", x"768f", x"768e", 
    x"768d", x"768c", x"768b", x"768a", x"7688", x"7687", x"7686", x"7685", 
    x"7684", x"7682", x"7681", x"7680", x"767f", x"767e", x"767d", x"767b", 
    x"767a", x"7679", x"7678", x"7677", x"7675", x"7674", x"7673", x"7672", 
    x"7671", x"766f", x"766e", x"766d", x"766c", x"766b", x"7669", x"7668", 
    x"7667", x"7666", x"7665", x"7664", x"7662", x"7661", x"7660", x"765f", 
    x"765e", x"765c", x"765b", x"765a", x"7659", x"7658", x"7656", x"7655", 
    x"7654", x"7653", x"7652", x"7650", x"764f", x"764e", x"764d", x"764c", 
    x"764a", x"7649", x"7648", x"7647", x"7646", x"7644", x"7643", x"7642", 
    x"7641", x"7640", x"763e", x"763d", x"763c", x"763b", x"763a", x"7638", 
    x"7637", x"7636", x"7635", x"7634", x"7632", x"7631", x"7630", x"762f", 
    x"762d", x"762c", x"762b", x"762a", x"7629", x"7627", x"7626", x"7625", 
    x"7624", x"7623", x"7621", x"7620", x"761f", x"761e", x"761d", x"761b", 
    x"761a", x"7619", x"7618", x"7617", x"7615", x"7614", x"7613", x"7612", 
    x"7610", x"760f", x"760e", x"760d", x"760c", x"760a", x"7609", x"7608", 
    x"7607", x"7606", x"7604", x"7603", x"7602", x"7601", x"75ff", x"75fe", 
    x"75fd", x"75fc", x"75fb", x"75f9", x"75f8", x"75f7", x"75f6", x"75f4", 
    x"75f3", x"75f2", x"75f1", x"75f0", x"75ee", x"75ed", x"75ec", x"75eb", 
    x"75e9", x"75e8", x"75e7", x"75e6", x"75e5", x"75e3", x"75e2", x"75e1", 
    x"75e0", x"75de", x"75dd", x"75dc", x"75db", x"75da", x"75d8", x"75d7", 
    x"75d6", x"75d5", x"75d3", x"75d2", x"75d1", x"75d0", x"75cf", x"75cd", 
    x"75cc", x"75cb", x"75ca", x"75c8", x"75c7", x"75c6", x"75c5", x"75c3", 
    x"75c2", x"75c1", x"75c0", x"75bf", x"75bd", x"75bc", x"75bb", x"75ba", 
    x"75b8", x"75b7", x"75b6", x"75b5", x"75b3", x"75b2", x"75b1", x"75b0", 
    x"75ae", x"75ad", x"75ac", x"75ab", x"75aa", x"75a8", x"75a7", x"75a6", 
    x"75a5", x"75a3", x"75a2", x"75a1", x"75a0", x"759e", x"759d", x"759c", 
    x"759b", x"7599", x"7598", x"7597", x"7596", x"7594", x"7593", x"7592", 
    x"7591", x"7590", x"758e", x"758d", x"758c", x"758b", x"7589", x"7588", 
    x"7587", x"7586", x"7584", x"7583", x"7582", x"7581", x"757f", x"757e", 
    x"757d", x"757c", x"757a", x"7579", x"7578", x"7577", x"7575", x"7574", 
    x"7573", x"7572", x"7570", x"756f", x"756e", x"756d", x"756b", x"756a", 
    x"7569", x"7568", x"7566", x"7565", x"7564", x"7563", x"7561", x"7560", 
    x"755f", x"755e", x"755c", x"755b", x"755a", x"7559", x"7557", x"7556", 
    x"7555", x"7554", x"7552", x"7551", x"7550", x"754f", x"754d", x"754c", 
    x"754b", x"754a", x"7548", x"7547", x"7546", x"7544", x"7543", x"7542", 
    x"7541", x"753f", x"753e", x"753d", x"753c", x"753a", x"7539", x"7538", 
    x"7537", x"7535", x"7534", x"7533", x"7532", x"7530", x"752f", x"752e", 
    x"752d", x"752b", x"752a", x"7529", x"7527", x"7526", x"7525", x"7524", 
    x"7522", x"7521", x"7520", x"751f", x"751d", x"751c", x"751b", x"751a", 
    x"7518", x"7517", x"7516", x"7514", x"7513", x"7512", x"7511", x"750f", 
    x"750e", x"750d", x"750c", x"750a", x"7509", x"7508", x"7506", x"7505", 
    x"7504", x"7503", x"7501", x"7500", x"74ff", x"74fe", x"74fc", x"74fb", 
    x"74fa", x"74f8", x"74f7", x"74f6", x"74f5", x"74f3", x"74f2", x"74f1", 
    x"74f0", x"74ee", x"74ed", x"74ec", x"74ea", x"74e9", x"74e8", x"74e7", 
    x"74e5", x"74e4", x"74e3", x"74e1", x"74e0", x"74df", x"74de", x"74dc", 
    x"74db", x"74da", x"74d8", x"74d7", x"74d6", x"74d5", x"74d3", x"74d2", 
    x"74d1", x"74cf", x"74ce", x"74cd", x"74cc", x"74ca", x"74c9", x"74c8", 
    x"74c6", x"74c5", x"74c4", x"74c3", x"74c1", x"74c0", x"74bf", x"74bd", 
    x"74bc", x"74bb", x"74ba", x"74b8", x"74b7", x"74b6", x"74b4", x"74b3", 
    x"74b2", x"74b1", x"74af", x"74ae", x"74ad", x"74ab", x"74aa", x"74a9", 
    x"74a8", x"74a6", x"74a5", x"74a4", x"74a2", x"74a1", x"74a0", x"749e", 
    x"749d", x"749c", x"749b", x"7499", x"7498", x"7497", x"7495", x"7494", 
    x"7493", x"7492", x"7490", x"748f", x"748e", x"748c", x"748b", x"748a", 
    x"7488", x"7487", x"7486", x"7485", x"7483", x"7482", x"7481", x"747f", 
    x"747e", x"747d", x"747b", x"747a", x"7479", x"7478", x"7476", x"7475", 
    x"7474", x"7472", x"7471", x"7470", x"746e", x"746d", x"746c", x"746a", 
    x"7469", x"7468", x"7467", x"7465", x"7464", x"7463", x"7461", x"7460", 
    x"745f", x"745d", x"745c", x"745b", x"7459", x"7458", x"7457", x"7456", 
    x"7454", x"7453", x"7452", x"7450", x"744f", x"744e", x"744c", x"744b", 
    x"744a", x"7448", x"7447", x"7446", x"7444", x"7443", x"7442", x"7441", 
    x"743f", x"743e", x"743d", x"743b", x"743a", x"7439", x"7437", x"7436", 
    x"7435", x"7433", x"7432", x"7431", x"742f", x"742e", x"742d", x"742b", 
    x"742a", x"7429", x"7428", x"7426", x"7425", x"7424", x"7422", x"7421", 
    x"7420", x"741e", x"741d", x"741c", x"741a", x"7419", x"7418", x"7416", 
    x"7415", x"7414", x"7412", x"7411", x"7410", x"740e", x"740d", x"740c", 
    x"740a", x"7409", x"7408", x"7406", x"7405", x"7404", x"7402", x"7401", 
    x"7400", x"73fe", x"73fd", x"73fc", x"73fa", x"73f9", x"73f8", x"73f7", 
    x"73f5", x"73f4", x"73f3", x"73f1", x"73f0", x"73ef", x"73ed", x"73ec", 
    x"73eb", x"73e9", x"73e8", x"73e7", x"73e5", x"73e4", x"73e3", x"73e1", 
    x"73e0", x"73df", x"73dd", x"73dc", x"73db", x"73d9", x"73d8", x"73d7", 
    x"73d5", x"73d4", x"73d3", x"73d1", x"73d0", x"73ce", x"73cd", x"73cc", 
    x"73ca", x"73c9", x"73c8", x"73c6", x"73c5", x"73c4", x"73c2", x"73c1", 
    x"73c0", x"73be", x"73bd", x"73bc", x"73ba", x"73b9", x"73b8", x"73b6", 
    x"73b5", x"73b4", x"73b2", x"73b1", x"73b0", x"73ae", x"73ad", x"73ac", 
    x"73aa", x"73a9", x"73a8", x"73a6", x"73a5", x"73a4", x"73a2", x"73a1", 
    x"739f", x"739e", x"739d", x"739b", x"739a", x"7399", x"7397", x"7396", 
    x"7395", x"7393", x"7392", x"7391", x"738f", x"738e", x"738d", x"738b", 
    x"738a", x"7389", x"7387", x"7386", x"7384", x"7383", x"7382", x"7380", 
    x"737f", x"737e", x"737c", x"737b", x"737a", x"7378", x"7377", x"7376", 
    x"7374", x"7373", x"7372", x"7370", x"736f", x"736d", x"736c", x"736b", 
    x"7369", x"7368", x"7367", x"7365", x"7364", x"7363", x"7361", x"7360", 
    x"735e", x"735d", x"735c", x"735a", x"7359", x"7358", x"7356", x"7355", 
    x"7354", x"7352", x"7351", x"7350", x"734e", x"734d", x"734b", x"734a", 
    x"7349", x"7347", x"7346", x"7345", x"7343", x"7342", x"7340", x"733f", 
    x"733e", x"733c", x"733b", x"733a", x"7338", x"7337", x"7336", x"7334", 
    x"7333", x"7331", x"7330", x"732f", x"732d", x"732c", x"732b", x"7329", 
    x"7328", x"7326", x"7325", x"7324", x"7322", x"7321", x"7320", x"731e", 
    x"731d", x"731c", x"731a", x"7319", x"7317", x"7316", x"7315", x"7313", 
    x"7312", x"7311", x"730f", x"730e", x"730c", x"730b", x"730a", x"7308", 
    x"7307", x"7305", x"7304", x"7303", x"7301", x"7300", x"72ff", x"72fd", 
    x"72fc", x"72fa", x"72f9", x"72f8", x"72f6", x"72f5", x"72f4", x"72f2", 
    x"72f1", x"72ef", x"72ee", x"72ed", x"72eb", x"72ea", x"72e8", x"72e7", 
    x"72e6", x"72e4", x"72e3", x"72e2", x"72e0", x"72df", x"72dd", x"72dc", 
    x"72db", x"72d9", x"72d8", x"72d6", x"72d5", x"72d4", x"72d2", x"72d1", 
    x"72d0", x"72ce", x"72cd", x"72cb", x"72ca", x"72c9", x"72c7", x"72c6", 
    x"72c4", x"72c3", x"72c2", x"72c0", x"72bf", x"72bd", x"72bc", x"72bb", 
    x"72b9", x"72b8", x"72b6", x"72b5", x"72b4", x"72b2", x"72b1", x"72b0", 
    x"72ae", x"72ad", x"72ab", x"72aa", x"72a9", x"72a7", x"72a6", x"72a4", 
    x"72a3", x"72a2", x"72a0", x"729f", x"729d", x"729c", x"729b", x"7299", 
    x"7298", x"7296", x"7295", x"7294", x"7292", x"7291", x"728f", x"728e", 
    x"728d", x"728b", x"728a", x"7288", x"7287", x"7286", x"7284", x"7283", 
    x"7281", x"7280", x"727f", x"727d", x"727c", x"727a", x"7279", x"7278", 
    x"7276", x"7275", x"7273", x"7272", x"7270", x"726f", x"726e", x"726c", 
    x"726b", x"7269", x"7268", x"7267", x"7265", x"7264", x"7262", x"7261", 
    x"7260", x"725e", x"725d", x"725b", x"725a", x"7259", x"7257", x"7256", 
    x"7254", x"7253", x"7251", x"7250", x"724f", x"724d", x"724c", x"724a", 
    x"7249", x"7248", x"7246", x"7245", x"7243", x"7242", x"7240", x"723f", 
    x"723e", x"723c", x"723b", x"7239", x"7238", x"7237", x"7235", x"7234", 
    x"7232", x"7231", x"722f", x"722e", x"722d", x"722b", x"722a", x"7228", 
    x"7227", x"7226", x"7224", x"7223", x"7221", x"7220", x"721e", x"721d", 
    x"721c", x"721a", x"7219", x"7217", x"7216", x"7214", x"7213", x"7212", 
    x"7210", x"720f", x"720d", x"720c", x"720a", x"7209", x"7208", x"7206", 
    x"7205", x"7203", x"7202", x"7200", x"71ff", x"71fe", x"71fc", x"71fb", 
    x"71f9", x"71f8", x"71f6", x"71f5", x"71f4", x"71f2", x"71f1", x"71ef", 
    x"71ee", x"71ec", x"71eb", x"71ea", x"71e8", x"71e7", x"71e5", x"71e4", 
    x"71e2", x"71e1", x"71e0", x"71de", x"71dd", x"71db", x"71da", x"71d8", 
    x"71d7", x"71d6", x"71d4", x"71d3", x"71d1", x"71d0", x"71ce", x"71cd", 
    x"71cb", x"71ca", x"71c9", x"71c7", x"71c6", x"71c4", x"71c3", x"71c1", 
    x"71c0", x"71be", x"71bd", x"71bc", x"71ba", x"71b9", x"71b7", x"71b6", 
    x"71b4", x"71b3", x"71b2", x"71b0", x"71af", x"71ad", x"71ac", x"71aa", 
    x"71a9", x"71a7", x"71a6", x"71a5", x"71a3", x"71a2", x"71a0", x"719f", 
    x"719d", x"719c", x"719a", x"7199", x"7197", x"7196", x"7195", x"7193", 
    x"7192", x"7190", x"718f", x"718d", x"718c", x"718a", x"7189", x"7188", 
    x"7186", x"7185", x"7183", x"7182", x"7180", x"717f", x"717d", x"717c", 
    x"717a", x"7179", x"7178", x"7176", x"7175", x"7173", x"7172", x"7170", 
    x"716f", x"716d", x"716c", x"716a", x"7169", x"7168", x"7166", x"7165", 
    x"7163", x"7162", x"7160", x"715f", x"715d", x"715c", x"715a", x"7159", 
    x"7158", x"7156", x"7155", x"7153", x"7152", x"7150", x"714f", x"714d", 
    x"714c", x"714a", x"7149", x"7147", x"7146", x"7145", x"7143", x"7142", 
    x"7140", x"713f", x"713d", x"713c", x"713a", x"7139", x"7137", x"7136", 
    x"7134", x"7133", x"7131", x"7130", x"712f", x"712d", x"712c", x"712a", 
    x"7129", x"7127", x"7126", x"7124", x"7123", x"7121", x"7120", x"711e", 
    x"711d", x"711b", x"711a", x"7119", x"7117", x"7116", x"7114", x"7113", 
    x"7111", x"7110", x"710e", x"710d", x"710b", x"710a", x"7108", x"7107", 
    x"7105", x"7104", x"7102", x"7101", x"70ff", x"70fe", x"70fd", x"70fb", 
    x"70fa", x"70f8", x"70f7", x"70f5", x"70f4", x"70f2", x"70f1", x"70ef", 
    x"70ee", x"70ec", x"70eb", x"70e9", x"70e8", x"70e6", x"70e5", x"70e3", 
    x"70e2", x"70e0", x"70df", x"70dd", x"70dc", x"70db", x"70d9", x"70d8", 
    x"70d6", x"70d5", x"70d3", x"70d2", x"70d0", x"70cf", x"70cd", x"70cc", 
    x"70ca", x"70c9", x"70c7", x"70c6", x"70c4", x"70c3", x"70c1", x"70c0", 
    x"70be", x"70bd", x"70bb", x"70ba", x"70b8", x"70b7", x"70b5", x"70b4", 
    x"70b2", x"70b1", x"70af", x"70ae", x"70ac", x"70ab", x"70a9", x"70a8", 
    x"70a6", x"70a5", x"70a3", x"70a2", x"70a0", x"709f", x"709e", x"709c", 
    x"709b", x"7099", x"7098", x"7096", x"7095", x"7093", x"7092", x"7090", 
    x"708f", x"708d", x"708c", x"708a", x"7089", x"7087", x"7086", x"7084", 
    x"7083", x"7081", x"7080", x"707e", x"707d", x"707b", x"707a", x"7078", 
    x"7077", x"7075", x"7074", x"7072", x"7071", x"706f", x"706e", x"706c", 
    x"706b", x"7069", x"7068", x"7066", x"7065", x"7063", x"7062", x"7060", 
    x"705f", x"705d", x"705c", x"705a", x"7059", x"7057", x"7056", x"7054", 
    x"7053", x"7051", x"7050", x"704e", x"704c", x"704b", x"7049", x"7048", 
    x"7046", x"7045", x"7043", x"7042", x"7040", x"703f", x"703d", x"703c", 
    x"703a", x"7039", x"7037", x"7036", x"7034", x"7033", x"7031", x"7030", 
    x"702e", x"702d", x"702b", x"702a", x"7028", x"7027", x"7025", x"7024", 
    x"7022", x"7021", x"701f", x"701e", x"701c", x"701b", x"7019", x"7018", 
    x"7016", x"7015", x"7013", x"7012", x"7010", x"700e", x"700d", x"700b", 
    x"700a", x"7008", x"7007", x"7005", x"7004", x"7002", x"7001", x"6fff", 
    x"6ffe", x"6ffc", x"6ffb", x"6ff9", x"6ff8", x"6ff6", x"6ff5", x"6ff3", 
    x"6ff2", x"6ff0", x"6fef", x"6fed", x"6feb", x"6fea", x"6fe8", x"6fe7", 
    x"6fe5", x"6fe4", x"6fe2", x"6fe1", x"6fdf", x"6fde", x"6fdc", x"6fdb", 
    x"6fd9", x"6fd8", x"6fd6", x"6fd5", x"6fd3", x"6fd2", x"6fd0", x"6fce", 
    x"6fcd", x"6fcb", x"6fca", x"6fc8", x"6fc7", x"6fc5", x"6fc4", x"6fc2", 
    x"6fc1", x"6fbf", x"6fbe", x"6fbc", x"6fbb", x"6fb9", x"6fb8", x"6fb6", 
    x"6fb4", x"6fb3", x"6fb1", x"6fb0", x"6fae", x"6fad", x"6fab", x"6faa", 
    x"6fa8", x"6fa7", x"6fa5", x"6fa4", x"6fa2", x"6fa0", x"6f9f", x"6f9d", 
    x"6f9c", x"6f9a", x"6f99", x"6f97", x"6f96", x"6f94", x"6f93", x"6f91", 
    x"6f90", x"6f8e", x"6f8c", x"6f8b", x"6f89", x"6f88", x"6f86", x"6f85", 
    x"6f83", x"6f82", x"6f80", x"6f7f", x"6f7d", x"6f7c", x"6f7a", x"6f78", 
    x"6f77", x"6f75", x"6f74", x"6f72", x"6f71", x"6f6f", x"6f6e", x"6f6c", 
    x"6f6b", x"6f69", x"6f67", x"6f66", x"6f64", x"6f63", x"6f61", x"6f60", 
    x"6f5e", x"6f5d", x"6f5b", x"6f59", x"6f58", x"6f56", x"6f55", x"6f53", 
    x"6f52", x"6f50", x"6f4f", x"6f4d", x"6f4c", x"6f4a", x"6f48", x"6f47", 
    x"6f45", x"6f44", x"6f42", x"6f41", x"6f3f", x"6f3e", x"6f3c", x"6f3a", 
    x"6f39", x"6f37", x"6f36", x"6f34", x"6f33", x"6f31", x"6f30", x"6f2e", 
    x"6f2c", x"6f2b", x"6f29", x"6f28", x"6f26", x"6f25", x"6f23", x"6f22", 
    x"6f20", x"6f1e", x"6f1d", x"6f1b", x"6f1a", x"6f18", x"6f17", x"6f15", 
    x"6f14", x"6f12", x"6f10", x"6f0f", x"6f0d", x"6f0c", x"6f0a", x"6f09", 
    x"6f07", x"6f05", x"6f04", x"6f02", x"6f01", x"6eff", x"6efe", x"6efc", 
    x"6efb", x"6ef9", x"6ef7", x"6ef6", x"6ef4", x"6ef3", x"6ef1", x"6ef0", 
    x"6eee", x"6eec", x"6eeb", x"6ee9", x"6ee8", x"6ee6", x"6ee5", x"6ee3", 
    x"6ee1", x"6ee0", x"6ede", x"6edd", x"6edb", x"6eda", x"6ed8", x"6ed6", 
    x"6ed5", x"6ed3", x"6ed2", x"6ed0", x"6ecf", x"6ecd", x"6ecb", x"6eca", 
    x"6ec8", x"6ec7", x"6ec5", x"6ec4", x"6ec2", x"6ec0", x"6ebf", x"6ebd", 
    x"6ebc", x"6eba", x"6eb9", x"6eb7", x"6eb5", x"6eb4", x"6eb2", x"6eb1", 
    x"6eaf", x"6ead", x"6eac", x"6eaa", x"6ea9", x"6ea7", x"6ea6", x"6ea4", 
    x"6ea2", x"6ea1", x"6e9f", x"6e9e", x"6e9c", x"6e9b", x"6e99", x"6e97", 
    x"6e96", x"6e94", x"6e93", x"6e91", x"6e8f", x"6e8e", x"6e8c", x"6e8b", 
    x"6e89", x"6e88", x"6e86", x"6e84", x"6e83", x"6e81", x"6e80", x"6e7e", 
    x"6e7c", x"6e7b", x"6e79", x"6e78", x"6e76", x"6e75", x"6e73", x"6e71", 
    x"6e70", x"6e6e", x"6e6d", x"6e6b", x"6e69", x"6e68", x"6e66", x"6e65", 
    x"6e63", x"6e61", x"6e60", x"6e5e", x"6e5d", x"6e5b", x"6e59", x"6e58", 
    x"6e56", x"6e55", x"6e53", x"6e52", x"6e50", x"6e4e", x"6e4d", x"6e4b", 
    x"6e4a", x"6e48", x"6e46", x"6e45", x"6e43", x"6e42", x"6e40", x"6e3e", 
    x"6e3d", x"6e3b", x"6e3a", x"6e38", x"6e36", x"6e35", x"6e33", x"6e32", 
    x"6e30", x"6e2e", x"6e2d", x"6e2b", x"6e2a", x"6e28", x"6e26", x"6e25", 
    x"6e23", x"6e22", x"6e20", x"6e1e", x"6e1d", x"6e1b", x"6e1a", x"6e18", 
    x"6e16", x"6e15", x"6e13", x"6e12", x"6e10", x"6e0e", x"6e0d", x"6e0b", 
    x"6e0a", x"6e08", x"6e06", x"6e05", x"6e03", x"6e02", x"6e00", x"6dfe", 
    x"6dfd", x"6dfb", x"6dfa", x"6df8", x"6df6", x"6df5", x"6df3", x"6df1", 
    x"6df0", x"6dee", x"6ded", x"6deb", x"6de9", x"6de8", x"6de6", x"6de5", 
    x"6de3", x"6de1", x"6de0", x"6dde", x"6ddd", x"6ddb", x"6dd9", x"6dd8", 
    x"6dd6", x"6dd4", x"6dd3", x"6dd1", x"6dd0", x"6dce", x"6dcc", x"6dcb", 
    x"6dc9", x"6dc8", x"6dc6", x"6dc4", x"6dc3", x"6dc1", x"6dbf", x"6dbe", 
    x"6dbc", x"6dbb", x"6db9", x"6db7", x"6db6", x"6db4", x"6db3", x"6db1", 
    x"6daf", x"6dae", x"6dac", x"6daa", x"6da9", x"6da7", x"6da6", x"6da4", 
    x"6da2", x"6da1", x"6d9f", x"6d9d", x"6d9c", x"6d9a", x"6d99", x"6d97", 
    x"6d95", x"6d94", x"6d92", x"6d91", x"6d8f", x"6d8d", x"6d8c", x"6d8a", 
    x"6d88", x"6d87", x"6d85", x"6d84", x"6d82", x"6d80", x"6d7f", x"6d7d", 
    x"6d7b", x"6d7a", x"6d78", x"6d76", x"6d75", x"6d73", x"6d72", x"6d70", 
    x"6d6e", x"6d6d", x"6d6b", x"6d69", x"6d68", x"6d66", x"6d65", x"6d63", 
    x"6d61", x"6d60", x"6d5e", x"6d5c", x"6d5b", x"6d59", x"6d58", x"6d56", 
    x"6d54", x"6d53", x"6d51", x"6d4f", x"6d4e", x"6d4c", x"6d4a", x"6d49", 
    x"6d47", x"6d46", x"6d44", x"6d42", x"6d41", x"6d3f", x"6d3d", x"6d3c", 
    x"6d3a", x"6d38", x"6d37", x"6d35", x"6d34", x"6d32", x"6d30", x"6d2f", 
    x"6d2d", x"6d2b", x"6d2a", x"6d28", x"6d26", x"6d25", x"6d23", x"6d21", 
    x"6d20", x"6d1e", x"6d1d", x"6d1b", x"6d19", x"6d18", x"6d16", x"6d14", 
    x"6d13", x"6d11", x"6d0f", x"6d0e", x"6d0c", x"6d0a", x"6d09", x"6d07", 
    x"6d06", x"6d04", x"6d02", x"6d01", x"6cff", x"6cfd", x"6cfc", x"6cfa", 
    x"6cf8", x"6cf7", x"6cf5", x"6cf3", x"6cf2", x"6cf0", x"6cee", x"6ced", 
    x"6ceb", x"6cea", x"6ce8", x"6ce6", x"6ce5", x"6ce3", x"6ce1", x"6ce0", 
    x"6cde", x"6cdc", x"6cdb", x"6cd9", x"6cd7", x"6cd6", x"6cd4", x"6cd2", 
    x"6cd1", x"6ccf", x"6ccd", x"6ccc", x"6cca", x"6cc8", x"6cc7", x"6cc5", 
    x"6cc3", x"6cc2", x"6cc0", x"6cbf", x"6cbd", x"6cbb", x"6cba", x"6cb8", 
    x"6cb6", x"6cb5", x"6cb3", x"6cb1", x"6cb0", x"6cae", x"6cac", x"6cab", 
    x"6ca9", x"6ca7", x"6ca6", x"6ca4", x"6ca2", x"6ca1", x"6c9f", x"6c9d", 
    x"6c9c", x"6c9a", x"6c98", x"6c97", x"6c95", x"6c93", x"6c92", x"6c90", 
    x"6c8e", x"6c8d", x"6c8b", x"6c89", x"6c88", x"6c86", x"6c84", x"6c83", 
    x"6c81", x"6c7f", x"6c7e", x"6c7c", x"6c7a", x"6c79", x"6c77", x"6c75", 
    x"6c74", x"6c72", x"6c70", x"6c6f", x"6c6d", x"6c6b", x"6c6a", x"6c68", 
    x"6c66", x"6c65", x"6c63", x"6c61", x"6c60", x"6c5e", x"6c5c", x"6c5b", 
    x"6c59", x"6c57", x"6c56", x"6c54", x"6c52", x"6c51", x"6c4f", x"6c4d", 
    x"6c4c", x"6c4a", x"6c48", x"6c47", x"6c45", x"6c43", x"6c42", x"6c40", 
    x"6c3e", x"6c3c", x"6c3b", x"6c39", x"6c37", x"6c36", x"6c34", x"6c32", 
    x"6c31", x"6c2f", x"6c2d", x"6c2c", x"6c2a", x"6c28", x"6c27", x"6c25", 
    x"6c23", x"6c22", x"6c20", x"6c1e", x"6c1d", x"6c1b", x"6c19", x"6c18", 
    x"6c16", x"6c14", x"6c12", x"6c11", x"6c0f", x"6c0d", x"6c0c", x"6c0a", 
    x"6c08", x"6c07", x"6c05", x"6c03", x"6c02", x"6c00", x"6bfe", x"6bfd", 
    x"6bfb", x"6bf9", x"6bf8", x"6bf6", x"6bf4", x"6bf2", x"6bf1", x"6bef", 
    x"6bed", x"6bec", x"6bea", x"6be8", x"6be7", x"6be5", x"6be3", x"6be2", 
    x"6be0", x"6bde", x"6bdd", x"6bdb", x"6bd9", x"6bd7", x"6bd6", x"6bd4", 
    x"6bd2", x"6bd1", x"6bcf", x"6bcd", x"6bcc", x"6bca", x"6bc8", x"6bc6", 
    x"6bc5", x"6bc3", x"6bc1", x"6bc0", x"6bbe", x"6bbc", x"6bbb", x"6bb9", 
    x"6bb7", x"6bb6", x"6bb4", x"6bb2", x"6bb0", x"6baf", x"6bad", x"6bab", 
    x"6baa", x"6ba8", x"6ba6", x"6ba5", x"6ba3", x"6ba1", x"6b9f", x"6b9e", 
    x"6b9c", x"6b9a", x"6b99", x"6b97", x"6b95", x"6b94", x"6b92", x"6b90", 
    x"6b8e", x"6b8d", x"6b8b", x"6b89", x"6b88", x"6b86", x"6b84", x"6b83", 
    x"6b81", x"6b7f", x"6b7d", x"6b7c", x"6b7a", x"6b78", x"6b77", x"6b75", 
    x"6b73", x"6b71", x"6b70", x"6b6e", x"6b6c", x"6b6b", x"6b69", x"6b67", 
    x"6b65", x"6b64", x"6b62", x"6b60", x"6b5f", x"6b5d", x"6b5b", x"6b5a", 
    x"6b58", x"6b56", x"6b54", x"6b53", x"6b51", x"6b4f", x"6b4e", x"6b4c", 
    x"6b4a", x"6b48", x"6b47", x"6b45", x"6b43", x"6b42", x"6b40", x"6b3e", 
    x"6b3c", x"6b3b", x"6b39", x"6b37", x"6b36", x"6b34", x"6b32", x"6b30", 
    x"6b2f", x"6b2d", x"6b2b", x"6b2a", x"6b28", x"6b26", x"6b24", x"6b23", 
    x"6b21", x"6b1f", x"6b1d", x"6b1c", x"6b1a", x"6b18", x"6b17", x"6b15", 
    x"6b13", x"6b11", x"6b10", x"6b0e", x"6b0c", x"6b0b", x"6b09", x"6b07", 
    x"6b05", x"6b04", x"6b02", x"6b00", x"6afe", x"6afd", x"6afb", x"6af9", 
    x"6af8", x"6af6", x"6af4", x"6af2", x"6af1", x"6aef", x"6aed", x"6aec", 
    x"6aea", x"6ae8", x"6ae6", x"6ae5", x"6ae3", x"6ae1", x"6adf", x"6ade", 
    x"6adc", x"6ada", x"6ad8", x"6ad7", x"6ad5", x"6ad3", x"6ad2", x"6ad0", 
    x"6ace", x"6acc", x"6acb", x"6ac9", x"6ac7", x"6ac5", x"6ac4", x"6ac2", 
    x"6ac0", x"6abf", x"6abd", x"6abb", x"6ab9", x"6ab8", x"6ab6", x"6ab4", 
    x"6ab2", x"6ab1", x"6aaf", x"6aad", x"6aab", x"6aaa", x"6aa8", x"6aa6", 
    x"6aa4", x"6aa3", x"6aa1", x"6a9f", x"6a9e", x"6a9c", x"6a9a", x"6a98", 
    x"6a97", x"6a95", x"6a93", x"6a91", x"6a90", x"6a8e", x"6a8c", x"6a8a", 
    x"6a89", x"6a87", x"6a85", x"6a83", x"6a82", x"6a80", x"6a7e", x"6a7c", 
    x"6a7b", x"6a79", x"6a77", x"6a75", x"6a74", x"6a72", x"6a70", x"6a6f", 
    x"6a6d", x"6a6b", x"6a69", x"6a68", x"6a66", x"6a64", x"6a62", x"6a61", 
    x"6a5f", x"6a5d", x"6a5b", x"6a5a", x"6a58", x"6a56", x"6a54", x"6a53", 
    x"6a51", x"6a4f", x"6a4d", x"6a4c", x"6a4a", x"6a48", x"6a46", x"6a45", 
    x"6a43", x"6a41", x"6a3f", x"6a3e", x"6a3c", x"6a3a", x"6a38", x"6a37", 
    x"6a35", x"6a33", x"6a31", x"6a30", x"6a2e", x"6a2c", x"6a2a", x"6a29", 
    x"6a27", x"6a25", x"6a23", x"6a21", x"6a20", x"6a1e", x"6a1c", x"6a1a", 
    x"6a19", x"6a17", x"6a15", x"6a13", x"6a12", x"6a10", x"6a0e", x"6a0c", 
    x"6a0b", x"6a09", x"6a07", x"6a05", x"6a04", x"6a02", x"6a00", x"69fe", 
    x"69fd", x"69fb", x"69f9", x"69f7", x"69f6", x"69f4", x"69f2", x"69f0", 
    x"69ee", x"69ed", x"69eb", x"69e9", x"69e7", x"69e6", x"69e4", x"69e2", 
    x"69e0", x"69df", x"69dd", x"69db", x"69d9", x"69d8", x"69d6", x"69d4", 
    x"69d2", x"69d0", x"69cf", x"69cd", x"69cb", x"69c9", x"69c8", x"69c6", 
    x"69c4", x"69c2", x"69c1", x"69bf", x"69bd", x"69bb", x"69b9", x"69b8", 
    x"69b6", x"69b4", x"69b2", x"69b1", x"69af", x"69ad", x"69ab", x"69a9", 
    x"69a8", x"69a6", x"69a4", x"69a2", x"69a1", x"699f", x"699d", x"699b", 
    x"699a", x"6998", x"6996", x"6994", x"6992", x"6991", x"698f", x"698d", 
    x"698b", x"698a", x"6988", x"6986", x"6984", x"6982", x"6981", x"697f", 
    x"697d", x"697b", x"697a", x"6978", x"6976", x"6974", x"6972", x"6971", 
    x"696f", x"696d", x"696b", x"696a", x"6968", x"6966", x"6964", x"6962", 
    x"6961", x"695f", x"695d", x"695b", x"6959", x"6958", x"6956", x"6954", 
    x"6952", x"6951", x"694f", x"694d", x"694b", x"6949", x"6948", x"6946", 
    x"6944", x"6942", x"6940", x"693f", x"693d", x"693b", x"6939", x"6938", 
    x"6936", x"6934", x"6932", x"6930", x"692f", x"692d", x"692b", x"6929", 
    x"6927", x"6926", x"6924", x"6922", x"6920", x"691e", x"691d", x"691b", 
    x"6919", x"6917", x"6915", x"6914", x"6912", x"6910", x"690e", x"690d", 
    x"690b", x"6909", x"6907", x"6905", x"6904", x"6902", x"6900", x"68fe", 
    x"68fc", x"68fb", x"68f9", x"68f7", x"68f5", x"68f3", x"68f2", x"68f0", 
    x"68ee", x"68ec", x"68ea", x"68e9", x"68e7", x"68e5", x"68e3", x"68e1", 
    x"68e0", x"68de", x"68dc", x"68da", x"68d8", x"68d7", x"68d5", x"68d3", 
    x"68d1", x"68cf", x"68ce", x"68cc", x"68ca", x"68c8", x"68c6", x"68c5", 
    x"68c3", x"68c1", x"68bf", x"68bd", x"68bb", x"68ba", x"68b8", x"68b6", 
    x"68b4", x"68b2", x"68b1", x"68af", x"68ad", x"68ab", x"68a9", x"68a8", 
    x"68a6", x"68a4", x"68a2", x"68a0", x"689f", x"689d", x"689b", x"6899", 
    x"6897", x"6896", x"6894", x"6892", x"6890", x"688e", x"688c", x"688b", 
    x"6889", x"6887", x"6885", x"6883", x"6882", x"6880", x"687e", x"687c", 
    x"687a", x"6879", x"6877", x"6875", x"6873", x"6871", x"686f", x"686e", 
    x"686c", x"686a", x"6868", x"6866", x"6865", x"6863", x"6861", x"685f", 
    x"685d", x"685b", x"685a", x"6858", x"6856", x"6854", x"6852", x"6851", 
    x"684f", x"684d", x"684b", x"6849", x"6847", x"6846", x"6844", x"6842", 
    x"6840", x"683e", x"683c", x"683b", x"6839", x"6837", x"6835", x"6833", 
    x"6832", x"6830", x"682e", x"682c", x"682a", x"6828", x"6827", x"6825", 
    x"6823", x"6821", x"681f", x"681d", x"681c", x"681a", x"6818", x"6816", 
    x"6814", x"6812", x"6811", x"680f", x"680d", x"680b", x"6809", x"6807", 
    x"6806", x"6804", x"6802", x"6800", x"67fe", x"67fd", x"67fb", x"67f9", 
    x"67f7", x"67f5", x"67f3", x"67f2", x"67f0", x"67ee", x"67ec", x"67ea", 
    x"67e8", x"67e7", x"67e5", x"67e3", x"67e1", x"67df", x"67dd", x"67dc", 
    x"67da", x"67d8", x"67d6", x"67d4", x"67d2", x"67d0", x"67cf", x"67cd", 
    x"67cb", x"67c9", x"67c7", x"67c5", x"67c4", x"67c2", x"67c0", x"67be", 
    x"67bc", x"67ba", x"67b9", x"67b7", x"67b5", x"67b3", x"67b1", x"67af", 
    x"67ae", x"67ac", x"67aa", x"67a8", x"67a6", x"67a4", x"67a2", x"67a1", 
    x"679f", x"679d", x"679b", x"6799", x"6797", x"6796", x"6794", x"6792", 
    x"6790", x"678e", x"678c", x"678a", x"6789", x"6787", x"6785", x"6783", 
    x"6781", x"677f", x"677e", x"677c", x"677a", x"6778", x"6776", x"6774", 
    x"6772", x"6771", x"676f", x"676d", x"676b", x"6769", x"6767", x"6765", 
    x"6764", x"6762", x"6760", x"675e", x"675c", x"675a", x"6759", x"6757", 
    x"6755", x"6753", x"6751", x"674f", x"674d", x"674c", x"674a", x"6748", 
    x"6746", x"6744", x"6742", x"6740", x"673f", x"673d", x"673b", x"6739", 
    x"6737", x"6735", x"6733", x"6732", x"6730", x"672e", x"672c", x"672a", 
    x"6728", x"6726", x"6725", x"6723", x"6721", x"671f", x"671d", x"671b", 
    x"6719", x"6718", x"6716", x"6714", x"6712", x"6710", x"670e", x"670c", 
    x"670a", x"6709", x"6707", x"6705", x"6703", x"6701", x"66ff", x"66fd", 
    x"66fc", x"66fa", x"66f8", x"66f6", x"66f4", x"66f2", x"66f0", x"66ee", 
    x"66ed", x"66eb", x"66e9", x"66e7", x"66e5", x"66e3", x"66e1", x"66e0", 
    x"66de", x"66dc", x"66da", x"66d8", x"66d6", x"66d4", x"66d2", x"66d1", 
    x"66cf", x"66cd", x"66cb", x"66c9", x"66c7", x"66c5", x"66c3", x"66c2", 
    x"66c0", x"66be", x"66bc", x"66ba", x"66b8", x"66b6", x"66b4", x"66b3", 
    x"66b1", x"66af", x"66ad", x"66ab", x"66a9", x"66a7", x"66a5", x"66a4", 
    x"66a2", x"66a0", x"669e", x"669c", x"669a", x"6698", x"6696", x"6695", 
    x"6693", x"6691", x"668f", x"668d", x"668b", x"6689", x"6687", x"6686", 
    x"6684", x"6682", x"6680", x"667e", x"667c", x"667a", x"6678", x"6676", 
    x"6675", x"6673", x"6671", x"666f", x"666d", x"666b", x"6669", x"6667", 
    x"6666", x"6664", x"6662", x"6660", x"665e", x"665c", x"665a", x"6658", 
    x"6656", x"6655", x"6653", x"6651", x"664f", x"664d", x"664b", x"6649", 
    x"6647", x"6645", x"6644", x"6642", x"6640", x"663e", x"663c", x"663a", 
    x"6638", x"6636", x"6634", x"6633", x"6631", x"662f", x"662d", x"662b", 
    x"6629", x"6627", x"6625", x"6623", x"6622", x"6620", x"661e", x"661c", 
    x"661a", x"6618", x"6616", x"6614", x"6612", x"6610", x"660f", x"660d", 
    x"660b", x"6609", x"6607", x"6605", x"6603", x"6601", x"65ff", x"65fd", 
    x"65fc", x"65fa", x"65f8", x"65f6", x"65f4", x"65f2", x"65f0", x"65ee", 
    x"65ec", x"65ea", x"65e9", x"65e7", x"65e5", x"65e3", x"65e1", x"65df", 
    x"65dd", x"65db", x"65d9", x"65d7", x"65d6", x"65d4", x"65d2", x"65d0", 
    x"65ce", x"65cc", x"65ca", x"65c8", x"65c6", x"65c4", x"65c3", x"65c1", 
    x"65bf", x"65bd", x"65bb", x"65b9", x"65b7", x"65b5", x"65b3", x"65b1", 
    x"65af", x"65ae", x"65ac", x"65aa", x"65a8", x"65a6", x"65a4", x"65a2", 
    x"65a0", x"659e", x"659c", x"659a", x"6599", x"6597", x"6595", x"6593", 
    x"6591", x"658f", x"658d", x"658b", x"6589", x"6587", x"6585", x"6584", 
    x"6582", x"6580", x"657e", x"657c", x"657a", x"6578", x"6576", x"6574", 
    x"6572", x"6570", x"656e", x"656d", x"656b", x"6569", x"6567", x"6565", 
    x"6563", x"6561", x"655f", x"655d", x"655b", x"6559", x"6557", x"6556", 
    x"6554", x"6552", x"6550", x"654e", x"654c", x"654a", x"6548", x"6546", 
    x"6544", x"6542", x"6540", x"653e", x"653d", x"653b", x"6539", x"6537", 
    x"6535", x"6533", x"6531", x"652f", x"652d", x"652b", x"6529", x"6527", 
    x"6525", x"6524", x"6522", x"6520", x"651e", x"651c", x"651a", x"6518", 
    x"6516", x"6514", x"6512", x"6510", x"650e", x"650c", x"650a", x"6509", 
    x"6507", x"6505", x"6503", x"6501", x"64ff", x"64fd", x"64fb", x"64f9", 
    x"64f7", x"64f5", x"64f3", x"64f1", x"64ef", x"64ee", x"64ec", x"64ea", 
    x"64e8", x"64e6", x"64e4", x"64e2", x"64e0", x"64de", x"64dc", x"64da", 
    x"64d8", x"64d6", x"64d4", x"64d2", x"64d1", x"64cf", x"64cd", x"64cb", 
    x"64c9", x"64c7", x"64c5", x"64c3", x"64c1", x"64bf", x"64bd", x"64bb", 
    x"64b9", x"64b7", x"64b5", x"64b3", x"64b2", x"64b0", x"64ae", x"64ac", 
    x"64aa", x"64a8", x"64a6", x"64a4", x"64a2", x"64a0", x"649e", x"649c", 
    x"649a", x"6498", x"6496", x"6494", x"6492", x"6491", x"648f", x"648d", 
    x"648b", x"6489", x"6487", x"6485", x"6483", x"6481", x"647f", x"647d", 
    x"647b", x"6479", x"6477", x"6475", x"6473", x"6471", x"646f", x"646e", 
    x"646c", x"646a", x"6468", x"6466", x"6464", x"6462", x"6460", x"645e", 
    x"645c", x"645a", x"6458", x"6456", x"6454", x"6452", x"6450", x"644e", 
    x"644c", x"644a", x"6448", x"6447", x"6445", x"6443", x"6441", x"643f", 
    x"643d", x"643b", x"6439", x"6437", x"6435", x"6433", x"6431", x"642f", 
    x"642d", x"642b", x"6429", x"6427", x"6425", x"6423", x"6421", x"641f", 
    x"641d", x"641c", x"641a", x"6418", x"6416", x"6414", x"6412", x"6410", 
    x"640e", x"640c", x"640a", x"6408", x"6406", x"6404", x"6402", x"6400", 
    x"63fe", x"63fc", x"63fa", x"63f8", x"63f6", x"63f4", x"63f2", x"63f0", 
    x"63ee", x"63ec", x"63ea", x"63e9", x"63e7", x"63e5", x"63e3", x"63e1", 
    x"63df", x"63dd", x"63db", x"63d9", x"63d7", x"63d5", x"63d3", x"63d1", 
    x"63cf", x"63cd", x"63cb", x"63c9", x"63c7", x"63c5", x"63c3", x"63c1", 
    x"63bf", x"63bd", x"63bb", x"63b9", x"63b7", x"63b5", x"63b3", x"63b1", 
    x"63af", x"63ae", x"63ac", x"63aa", x"63a8", x"63a6", x"63a4", x"63a2", 
    x"63a0", x"639e", x"639c", x"639a", x"6398", x"6396", x"6394", x"6392", 
    x"6390", x"638e", x"638c", x"638a", x"6388", x"6386", x"6384", x"6382", 
    x"6380", x"637e", x"637c", x"637a", x"6378", x"6376", x"6374", x"6372", 
    x"6370", x"636e", x"636c", x"636a", x"6368", x"6366", x"6364", x"6362", 
    x"6360", x"635e", x"635d", x"635b", x"6359", x"6357", x"6355", x"6353", 
    x"6351", x"634f", x"634d", x"634b", x"6349", x"6347", x"6345", x"6343", 
    x"6341", x"633f", x"633d", x"633b", x"6339", x"6337", x"6335", x"6333", 
    x"6331", x"632f", x"632d", x"632b", x"6329", x"6327", x"6325", x"6323", 
    x"6321", x"631f", x"631d", x"631b", x"6319", x"6317", x"6315", x"6313", 
    x"6311", x"630f", x"630d", x"630b", x"6309", x"6307", x"6305", x"6303", 
    x"6301", x"62ff", x"62fd", x"62fb", x"62f9", x"62f7", x"62f5", x"62f3", 
    x"62f1", x"62ef", x"62ed", x"62eb", x"62e9", x"62e7", x"62e5", x"62e3", 
    x"62e1", x"62df", x"62dd", x"62db", x"62d9", x"62d7", x"62d5", x"62d3", 
    x"62d1", x"62cf", x"62cd", x"62cb", x"62c9", x"62c7", x"62c5", x"62c3", 
    x"62c1", x"62bf", x"62bd", x"62bb", x"62b9", x"62b7", x"62b5", x"62b3", 
    x"62b1", x"62af", x"62ad", x"62ab", x"62a9", x"62a7", x"62a5", x"62a3", 
    x"62a1", x"629f", x"629d", x"629b", x"6299", x"6297", x"6295", x"6293", 
    x"6291", x"628f", x"628d", x"628b", x"6289", x"6287", x"6285", x"6283", 
    x"6281", x"627f", x"627d", x"627b", x"6279", x"6277", x"6275", x"6273", 
    x"6271", x"626f", x"626d", x"626b", x"6269", x"6267", x"6265", x"6263", 
    x"6261", x"625f", x"625d", x"625b", x"6259", x"6257", x"6255", x"6253", 
    x"6251", x"624f", x"624d", x"624b", x"6249", x"6247", x"6245", x"6243", 
    x"6241", x"623f", x"623d", x"623b", x"6239", x"6237", x"6235", x"6233", 
    x"6231", x"622f", x"622d", x"622b", x"6229", x"6227", x"6225", x"6223", 
    x"6221", x"621f", x"621d", x"621b", x"6219", x"6217", x"6215", x"6213", 
    x"6211", x"620f", x"620d", x"620b", x"6208", x"6206", x"6204", x"6202", 
    x"6200", x"61fe", x"61fc", x"61fa", x"61f8", x"61f6", x"61f4", x"61f2", 
    x"61f0", x"61ee", x"61ec", x"61ea", x"61e8", x"61e6", x"61e4", x"61e2", 
    x"61e0", x"61de", x"61dc", x"61da", x"61d8", x"61d6", x"61d4", x"61d2", 
    x"61d0", x"61ce", x"61cc", x"61ca", x"61c8", x"61c6", x"61c4", x"61c2", 
    x"61c0", x"61be", x"61bc", x"61ba", x"61b8", x"61b5", x"61b3", x"61b1", 
    x"61af", x"61ad", x"61ab", x"61a9", x"61a7", x"61a5", x"61a3", x"61a1", 
    x"619f", x"619d", x"619b", x"6199", x"6197", x"6195", x"6193", x"6191", 
    x"618f", x"618d", x"618b", x"6189", x"6187", x"6185", x"6183", x"6181", 
    x"617f", x"617d", x"617b", x"6179", x"6176", x"6174", x"6172", x"6170", 
    x"616e", x"616c", x"616a", x"6168", x"6166", x"6164", x"6162", x"6160", 
    x"615e", x"615c", x"615a", x"6158", x"6156", x"6154", x"6152", x"6150", 
    x"614e", x"614c", x"614a", x"6148", x"6146", x"6143", x"6141", x"613f", 
    x"613d", x"613b", x"6139", x"6137", x"6135", x"6133", x"6131", x"612f", 
    x"612d", x"612b", x"6129", x"6127", x"6125", x"6123", x"6121", x"611f", 
    x"611d", x"611b", x"6119", x"6117", x"6114", x"6112", x"6110", x"610e", 
    x"610c", x"610a", x"6108", x"6106", x"6104", x"6102", x"6100", x"60fe", 
    x"60fc", x"60fa", x"60f8", x"60f6", x"60f4", x"60f2", x"60f0", x"60ee", 
    x"60eb", x"60e9", x"60e7", x"60e5", x"60e3", x"60e1", x"60df", x"60dd", 
    x"60db", x"60d9", x"60d7", x"60d5", x"60d3", x"60d1", x"60cf", x"60cd", 
    x"60cb", x"60c9", x"60c6", x"60c4", x"60c2", x"60c0", x"60be", x"60bc", 
    x"60ba", x"60b8", x"60b6", x"60b4", x"60b2", x"60b0", x"60ae", x"60ac", 
    x"60aa", x"60a8", x"60a6", x"60a4", x"60a1", x"609f", x"609d", x"609b", 
    x"6099", x"6097", x"6095", x"6093", x"6091", x"608f", x"608d", x"608b", 
    x"6089", x"6087", x"6085", x"6083", x"6080", x"607e", x"607c", x"607a", 
    x"6078", x"6076", x"6074", x"6072", x"6070", x"606e", x"606c", x"606a", 
    x"6068", x"6066", x"6064", x"6061", x"605f", x"605d", x"605b", x"6059", 
    x"6057", x"6055", x"6053", x"6051", x"604f", x"604d", x"604b", x"6049", 
    x"6047", x"6045", x"6042", x"6040", x"603e", x"603c", x"603a", x"6038", 
    x"6036", x"6034", x"6032", x"6030", x"602e", x"602c", x"602a", x"6028", 
    x"6025", x"6023", x"6021", x"601f", x"601d", x"601b", x"6019", x"6017", 
    x"6015", x"6013", x"6011", x"600f", x"600d", x"600a", x"6008", x"6006", 
    x"6004", x"6002", x"6000", x"5ffe", x"5ffc", x"5ffa", x"5ff8", x"5ff6", 
    x"5ff4", x"5ff2", x"5fef", x"5fed", x"5feb", x"5fe9", x"5fe7", x"5fe5", 
    x"5fe3", x"5fe1", x"5fdf", x"5fdd", x"5fdb", x"5fd9", x"5fd6", x"5fd4", 
    x"5fd2", x"5fd0", x"5fce", x"5fcc", x"5fca", x"5fc8", x"5fc6", x"5fc4", 
    x"5fc2", x"5fc0", x"5fbd", x"5fbb", x"5fb9", x"5fb7", x"5fb5", x"5fb3", 
    x"5fb1", x"5faf", x"5fad", x"5fab", x"5fa9", x"5fa7", x"5fa4", x"5fa2", 
    x"5fa0", x"5f9e", x"5f9c", x"5f9a", x"5f98", x"5f96", x"5f94", x"5f92", 
    x"5f90", x"5f8d", x"5f8b", x"5f89", x"5f87", x"5f85", x"5f83", x"5f81", 
    x"5f7f", x"5f7d", x"5f7b", x"5f79", x"5f76", x"5f74", x"5f72", x"5f70", 
    x"5f6e", x"5f6c", x"5f6a", x"5f68", x"5f66", x"5f64", x"5f61", x"5f5f", 
    x"5f5d", x"5f5b", x"5f59", x"5f57", x"5f55", x"5f53", x"5f51", x"5f4f", 
    x"5f4d", x"5f4a", x"5f48", x"5f46", x"5f44", x"5f42", x"5f40", x"5f3e", 
    x"5f3c", x"5f3a", x"5f38", x"5f35", x"5f33", x"5f31", x"5f2f", x"5f2d", 
    x"5f2b", x"5f29", x"5f27", x"5f25", x"5f23", x"5f20", x"5f1e", x"5f1c", 
    x"5f1a", x"5f18", x"5f16", x"5f14", x"5f12", x"5f10", x"5f0e", x"5f0b", 
    x"5f09", x"5f07", x"5f05", x"5f03", x"5f01", x"5eff", x"5efd", x"5efb", 
    x"5ef8", x"5ef6", x"5ef4", x"5ef2", x"5ef0", x"5eee", x"5eec", x"5eea", 
    x"5ee8", x"5ee6", x"5ee3", x"5ee1", x"5edf", x"5edd", x"5edb", x"5ed9", 
    x"5ed7", x"5ed5", x"5ed3", x"5ed0", x"5ece", x"5ecc", x"5eca", x"5ec8", 
    x"5ec6", x"5ec4", x"5ec2", x"5ec0", x"5ebd", x"5ebb", x"5eb9", x"5eb7", 
    x"5eb5", x"5eb3", x"5eb1", x"5eaf", x"5ead", x"5eaa", x"5ea8", x"5ea6", 
    x"5ea4", x"5ea2", x"5ea0", x"5e9e", x"5e9c", x"5e99", x"5e97", x"5e95", 
    x"5e93", x"5e91", x"5e8f", x"5e8d", x"5e8b", x"5e89", x"5e86", x"5e84", 
    x"5e82", x"5e80", x"5e7e", x"5e7c", x"5e7a", x"5e78", x"5e75", x"5e73", 
    x"5e71", x"5e6f", x"5e6d", x"5e6b", x"5e69", x"5e67", x"5e64", x"5e62", 
    x"5e60", x"5e5e", x"5e5c", x"5e5a", x"5e58", x"5e56", x"5e54", x"5e51", 
    x"5e4f", x"5e4d", x"5e4b", x"5e49", x"5e47", x"5e45", x"5e43", x"5e40", 
    x"5e3e", x"5e3c", x"5e3a", x"5e38", x"5e36", x"5e34", x"5e32", x"5e2f", 
    x"5e2d", x"5e2b", x"5e29", x"5e27", x"5e25", x"5e23", x"5e20", x"5e1e", 
    x"5e1c", x"5e1a", x"5e18", x"5e16", x"5e14", x"5e12", x"5e0f", x"5e0d", 
    x"5e0b", x"5e09", x"5e07", x"5e05", x"5e03", x"5e01", x"5dfe", x"5dfc", 
    x"5dfa", x"5df8", x"5df6", x"5df4", x"5df2", x"5def", x"5ded", x"5deb", 
    x"5de9", x"5de7", x"5de5", x"5de3", x"5de1", x"5dde", x"5ddc", x"5dda", 
    x"5dd8", x"5dd6", x"5dd4", x"5dd2", x"5dcf", x"5dcd", x"5dcb", x"5dc9", 
    x"5dc7", x"5dc5", x"5dc3", x"5dc0", x"5dbe", x"5dbc", x"5dba", x"5db8", 
    x"5db6", x"5db4", x"5db1", x"5daf", x"5dad", x"5dab", x"5da9", x"5da7", 
    x"5da5", x"5da3", x"5da0", x"5d9e", x"5d9c", x"5d9a", x"5d98", x"5d96", 
    x"5d94", x"5d91", x"5d8f", x"5d8d", x"5d8b", x"5d89", x"5d87", x"5d84", 
    x"5d82", x"5d80", x"5d7e", x"5d7c", x"5d7a", x"5d78", x"5d75", x"5d73", 
    x"5d71", x"5d6f", x"5d6d", x"5d6b", x"5d69", x"5d66", x"5d64", x"5d62", 
    x"5d60", x"5d5e", x"5d5c", x"5d5a", x"5d57", x"5d55", x"5d53", x"5d51", 
    x"5d4f", x"5d4d", x"5d4b", x"5d48", x"5d46", x"5d44", x"5d42", x"5d40", 
    x"5d3e", x"5d3b", x"5d39", x"5d37", x"5d35", x"5d33", x"5d31", x"5d2f", 
    x"5d2c", x"5d2a", x"5d28", x"5d26", x"5d24", x"5d22", x"5d1f", x"5d1d", 
    x"5d1b", x"5d19", x"5d17", x"5d15", x"5d13", x"5d10", x"5d0e", x"5d0c", 
    x"5d0a", x"5d08", x"5d06", x"5d03", x"5d01", x"5cff", x"5cfd", x"5cfb", 
    x"5cf9", x"5cf6", x"5cf4", x"5cf2", x"5cf0", x"5cee", x"5cec", x"5ce9", 
    x"5ce7", x"5ce5", x"5ce3", x"5ce1", x"5cdf", x"5cdd", x"5cda", x"5cd8", 
    x"5cd6", x"5cd4", x"5cd2", x"5cd0", x"5ccd", x"5ccb", x"5cc9", x"5cc7", 
    x"5cc5", x"5cc3", x"5cc0", x"5cbe", x"5cbc", x"5cba", x"5cb8", x"5cb6", 
    x"5cb3", x"5cb1", x"5caf", x"5cad", x"5cab", x"5ca9", x"5ca6", x"5ca4", 
    x"5ca2", x"5ca0", x"5c9e", x"5c9c", x"5c99", x"5c97", x"5c95", x"5c93", 
    x"5c91", x"5c8f", x"5c8c", x"5c8a", x"5c88", x"5c86", x"5c84", x"5c82", 
    x"5c7f", x"5c7d", x"5c7b", x"5c79", x"5c77", x"5c74", x"5c72", x"5c70", 
    x"5c6e", x"5c6c", x"5c6a", x"5c67", x"5c65", x"5c63", x"5c61", x"5c5f", 
    x"5c5d", x"5c5a", x"5c58", x"5c56", x"5c54", x"5c52", x"5c50", x"5c4d", 
    x"5c4b", x"5c49", x"5c47", x"5c45", x"5c42", x"5c40", x"5c3e", x"5c3c", 
    x"5c3a", x"5c38", x"5c35", x"5c33", x"5c31", x"5c2f", x"5c2d", x"5c2b", 
    x"5c28", x"5c26", x"5c24", x"5c22", x"5c20", x"5c1d", x"5c1b", x"5c19", 
    x"5c17", x"5c15", x"5c13", x"5c10", x"5c0e", x"5c0c", x"5c0a", x"5c08", 
    x"5c05", x"5c03", x"5c01", x"5bff", x"5bfd", x"5bfa", x"5bf8", x"5bf6", 
    x"5bf4", x"5bf2", x"5bf0", x"5bed", x"5beb", x"5be9", x"5be7", x"5be5", 
    x"5be2", x"5be0", x"5bde", x"5bdc", x"5bda", x"5bd8", x"5bd5", x"5bd3", 
    x"5bd1", x"5bcf", x"5bcd", x"5bca", x"5bc8", x"5bc6", x"5bc4", x"5bc2", 
    x"5bbf", x"5bbd", x"5bbb", x"5bb9", x"5bb7", x"5bb4", x"5bb2", x"5bb0", 
    x"5bae", x"5bac", x"5baa", x"5ba7", x"5ba5", x"5ba3", x"5ba1", x"5b9f", 
    x"5b9c", x"5b9a", x"5b98", x"5b96", x"5b94", x"5b91", x"5b8f", x"5b8d", 
    x"5b8b", x"5b89", x"5b86", x"5b84", x"5b82", x"5b80", x"5b7e", x"5b7b", 
    x"5b79", x"5b77", x"5b75", x"5b73", x"5b70", x"5b6e", x"5b6c", x"5b6a", 
    x"5b68", x"5b65", x"5b63", x"5b61", x"5b5f", x"5b5d", x"5b5a", x"5b58", 
    x"5b56", x"5b54", x"5b52", x"5b4f", x"5b4d", x"5b4b", x"5b49", x"5b47", 
    x"5b44", x"5b42", x"5b40", x"5b3e", x"5b3c", x"5b39", x"5b37", x"5b35", 
    x"5b33", x"5b31", x"5b2e", x"5b2c", x"5b2a", x"5b28", x"5b26", x"5b23", 
    x"5b21", x"5b1f", x"5b1d", x"5b1b", x"5b18", x"5b16", x"5b14", x"5b12", 
    x"5b0f", x"5b0d", x"5b0b", x"5b09", x"5b07", x"5b04", x"5b02", x"5b00", 
    x"5afe", x"5afc", x"5af9", x"5af7", x"5af5", x"5af3", x"5af1", x"5aee", 
    x"5aec", x"5aea", x"5ae8", x"5ae6", x"5ae3", x"5ae1", x"5adf", x"5add", 
    x"5ada", x"5ad8", x"5ad6", x"5ad4", x"5ad2", x"5acf", x"5acd", x"5acb", 
    x"5ac9", x"5ac7", x"5ac4", x"5ac2", x"5ac0", x"5abe", x"5abb", x"5ab9", 
    x"5ab7", x"5ab5", x"5ab3", x"5ab0", x"5aae", x"5aac", x"5aaa", x"5aa8", 
    x"5aa5", x"5aa3", x"5aa1", x"5a9f", x"5a9c", x"5a9a", x"5a98", x"5a96", 
    x"5a94", x"5a91", x"5a8f", x"5a8d", x"5a8b", x"5a88", x"5a86", x"5a84", 
    x"5a82", x"5a80", x"5a7d", x"5a7b", x"5a79", x"5a77", x"5a74", x"5a72", 
    x"5a70", x"5a6e", x"5a6c", x"5a69", x"5a67", x"5a65", x"5a63", x"5a60", 
    x"5a5e", x"5a5c", x"5a5a", x"5a58", x"5a55", x"5a53", x"5a51", x"5a4f", 
    x"5a4c", x"5a4a", x"5a48", x"5a46", x"5a43", x"5a41", x"5a3f", x"5a3d", 
    x"5a3b", x"5a38", x"5a36", x"5a34", x"5a32", x"5a2f", x"5a2d", x"5a2b", 
    x"5a29", x"5a27", x"5a24", x"5a22", x"5a20", x"5a1e", x"5a1b", x"5a19", 
    x"5a17", x"5a15", x"5a12", x"5a10", x"5a0e", x"5a0c", x"5a0a", x"5a07", 
    x"5a05", x"5a03", x"5a01", x"59fe", x"59fc", x"59fa", x"59f8", x"59f5", 
    x"59f3", x"59f1", x"59ef", x"59ec", x"59ea", x"59e8", x"59e6", x"59e4", 
    x"59e1", x"59df", x"59dd", x"59db", x"59d8", x"59d6", x"59d4", x"59d2", 
    x"59cf", x"59cd", x"59cb", x"59c9", x"59c6", x"59c4", x"59c2", x"59c0", 
    x"59bd", x"59bb", x"59b9", x"59b7", x"59b5", x"59b2", x"59b0", x"59ae", 
    x"59ac", x"59a9", x"59a7", x"59a5", x"59a3", x"59a0", x"599e", x"599c", 
    x"599a", x"5997", x"5995", x"5993", x"5991", x"598e", x"598c", x"598a", 
    x"5988", x"5985", x"5983", x"5981", x"597f", x"597c", x"597a", x"5978", 
    x"5976", x"5973", x"5971", x"596f", x"596d", x"596a", x"5968", x"5966", 
    x"5964", x"5961", x"595f", x"595d", x"595b", x"5958", x"5956", x"5954", 
    x"5952", x"594f", x"594d", x"594b", x"5949", x"5946", x"5944", x"5942", 
    x"5940", x"593d", x"593b", x"5939", x"5937", x"5934", x"5932", x"5930", 
    x"592e", x"592b", x"5929", x"5927", x"5925", x"5922", x"5920", x"591e", 
    x"591c", x"5919", x"5917", x"5915", x"5913", x"5910", x"590e", x"590c", 
    x"590a", x"5907", x"5905", x"5903", x"5901", x"58fe", x"58fc", x"58fa", 
    x"58f8", x"58f5", x"58f3", x"58f1", x"58ee", x"58ec", x"58ea", x"58e8", 
    x"58e5", x"58e3", x"58e1", x"58df", x"58dc", x"58da", x"58d8", x"58d6", 
    x"58d3", x"58d1", x"58cf", x"58cd", x"58ca", x"58c8", x"58c6", x"58c4", 
    x"58c1", x"58bf", x"58bd", x"58ba", x"58b8", x"58b6", x"58b4", x"58b1", 
    x"58af", x"58ad", x"58ab", x"58a8", x"58a6", x"58a4", x"58a2", x"589f", 
    x"589d", x"589b", x"5898", x"5896", x"5894", x"5892", x"588f", x"588d", 
    x"588b", x"5889", x"5886", x"5884", x"5882", x"5880", x"587d", x"587b", 
    x"5879", x"5876", x"5874", x"5872", x"5870", x"586d", x"586b", x"5869", 
    x"5867", x"5864", x"5862", x"5860", x"585d", x"585b", x"5859", x"5857", 
    x"5854", x"5852", x"5850", x"584e", x"584b", x"5849", x"5847", x"5844", 
    x"5842", x"5840", x"583e", x"583b", x"5839", x"5837", x"5835", x"5832", 
    x"5830", x"582e", x"582b", x"5829", x"5827", x"5825", x"5822", x"5820", 
    x"581e", x"581b", x"5819", x"5817", x"5815", x"5812", x"5810", x"580e", 
    x"580c", x"5809", x"5807", x"5805", x"5802", x"5800", x"57fe", x"57fc", 
    x"57f9", x"57f7", x"57f5", x"57f2", x"57f0", x"57ee", x"57ec", x"57e9", 
    x"57e7", x"57e5", x"57e2", x"57e0", x"57de", x"57dc", x"57d9", x"57d7", 
    x"57d5", x"57d2", x"57d0", x"57ce", x"57cc", x"57c9", x"57c7", x"57c5", 
    x"57c2", x"57c0", x"57be", x"57bc", x"57b9", x"57b7", x"57b5", x"57b2", 
    x"57b0", x"57ae", x"57ac", x"57a9", x"57a7", x"57a5", x"57a2", x"57a0", 
    x"579e", x"579c", x"5799", x"5797", x"5795", x"5792", x"5790", x"578e", 
    x"578b", x"5789", x"5787", x"5785", x"5782", x"5780", x"577e", x"577b", 
    x"5779", x"5777", x"5775", x"5772", x"5770", x"576e", x"576b", x"5769", 
    x"5767", x"5765", x"5762", x"5760", x"575e", x"575b", x"5759", x"5757", 
    x"5754", x"5752", x"5750", x"574e", x"574b", x"5749", x"5747", x"5744", 
    x"5742", x"5740", x"573d", x"573b", x"5739", x"5737", x"5734", x"5732", 
    x"5730", x"572d", x"572b", x"5729", x"5726", x"5724", x"5722", x"5720", 
    x"571d", x"571b", x"5719", x"5716", x"5714", x"5712", x"570f", x"570d", 
    x"570b", x"5709", x"5706", x"5704", x"5702", x"56ff", x"56fd", x"56fb", 
    x"56f8", x"56f6", x"56f4", x"56f1", x"56ef", x"56ed", x"56eb", x"56e8", 
    x"56e6", x"56e4", x"56e1", x"56df", x"56dd", x"56da", x"56d8", x"56d6", 
    x"56d3", x"56d1", x"56cf", x"56cd", x"56ca", x"56c8", x"56c6", x"56c3", 
    x"56c1", x"56bf", x"56bc", x"56ba", x"56b8", x"56b5", x"56b3", x"56b1", 
    x"56af", x"56ac", x"56aa", x"56a8", x"56a5", x"56a3", x"56a1", x"569e", 
    x"569c", x"569a", x"5697", x"5695", x"5693", x"5690", x"568e", x"568c", 
    x"568a", x"5687", x"5685", x"5683", x"5680", x"567e", x"567c", x"5679", 
    x"5677", x"5675", x"5672", x"5670", x"566e", x"566b", x"5669", x"5667", 
    x"5664", x"5662", x"5660", x"565e", x"565b", x"5659", x"5657", x"5654", 
    x"5652", x"5650", x"564d", x"564b", x"5649", x"5646", x"5644", x"5642", 
    x"563f", x"563d", x"563b", x"5638", x"5636", x"5634", x"5631", x"562f", 
    x"562d", x"562a", x"5628", x"5626", x"5623", x"5621", x"561f", x"561d", 
    x"561a", x"5618", x"5616", x"5613", x"5611", x"560f", x"560c", x"560a", 
    x"5608", x"5605", x"5603", x"5601", x"55fe", x"55fc", x"55fa", x"55f7", 
    x"55f5", x"55f3", x"55f0", x"55ee", x"55ec", x"55e9", x"55e7", x"55e5", 
    x"55e2", x"55e0", x"55de", x"55db", x"55d9", x"55d7", x"55d4", x"55d2", 
    x"55d0", x"55cd", x"55cb", x"55c9", x"55c6", x"55c4", x"55c2", x"55bf", 
    x"55bd", x"55bb", x"55b8", x"55b6", x"55b4", x"55b1", x"55af", x"55ad", 
    x"55aa", x"55a8", x"55a6", x"55a3", x"55a1", x"559f", x"559c", x"559a", 
    x"5598", x"5595", x"5593", x"5591", x"558e", x"558c", x"558a", x"5587", 
    x"5585", x"5583", x"5580", x"557e", x"557c", x"5579", x"5577", x"5575", 
    x"5572", x"5570", x"556e", x"556b", x"5569", x"5567", x"5564", x"5562", 
    x"5560", x"555d", x"555b", x"5559", x"5556", x"5554", x"5552", x"554f", 
    x"554d", x"554b", x"5548", x"5546", x"5543", x"5541", x"553f", x"553c", 
    x"553a", x"5538", x"5535", x"5533", x"5531", x"552e", x"552c", x"552a", 
    x"5527", x"5525", x"5523", x"5520", x"551e", x"551c", x"5519", x"5517", 
    x"5515", x"5512", x"5510", x"550e", x"550b", x"5509", x"5506", x"5504", 
    x"5502", x"54ff", x"54fd", x"54fb", x"54f8", x"54f6", x"54f4", x"54f1", 
    x"54ef", x"54ed", x"54ea", x"54e8", x"54e6", x"54e3", x"54e1", x"54df", 
    x"54dc", x"54da", x"54d7", x"54d5", x"54d3", x"54d0", x"54ce", x"54cc", 
    x"54c9", x"54c7", x"54c5", x"54c2", x"54c0", x"54be", x"54bb", x"54b9", 
    x"54b7", x"54b4", x"54b2", x"54af", x"54ad", x"54ab", x"54a8", x"54a6", 
    x"54a4", x"54a1", x"549f", x"549d", x"549a", x"5498", x"5496", x"5493", 
    x"5491", x"548e", x"548c", x"548a", x"5487", x"5485", x"5483", x"5480", 
    x"547e", x"547c", x"5479", x"5477", x"5475", x"5472", x"5470", x"546d", 
    x"546b", x"5469", x"5466", x"5464", x"5462", x"545f", x"545d", x"545b", 
    x"5458", x"5456", x"5453", x"5451", x"544f", x"544c", x"544a", x"5448", 
    x"5445", x"5443", x"5441", x"543e", x"543c", x"5439", x"5437", x"5435", 
    x"5432", x"5430", x"542e", x"542b", x"5429", x"5427", x"5424", x"5422", 
    x"541f", x"541d", x"541b", x"5418", x"5416", x"5414", x"5411", x"540f", 
    x"540c", x"540a", x"5408", x"5405", x"5403", x"5401", x"53fe", x"53fc", 
    x"53fa", x"53f7", x"53f5", x"53f2", x"53f0", x"53ee", x"53eb", x"53e9", 
    x"53e7", x"53e4", x"53e2", x"53df", x"53dd", x"53db", x"53d8", x"53d6", 
    x"53d4", x"53d1", x"53cf", x"53cc", x"53ca", x"53c8", x"53c5", x"53c3", 
    x"53c1", x"53be", x"53bc", x"53b9", x"53b7", x"53b5", x"53b2", x"53b0", 
    x"53ae", x"53ab", x"53a9", x"53a6", x"53a4", x"53a2", x"539f", x"539d", 
    x"539b", x"5398", x"5396", x"5393", x"5391", x"538f", x"538c", x"538a", 
    x"5387", x"5385", x"5383", x"5380", x"537e", x"537c", x"5379", x"5377", 
    x"5374", x"5372", x"5370", x"536d", x"536b", x"5369", x"5366", x"5364", 
    x"5361", x"535f", x"535d", x"535a", x"5358", x"5355", x"5353", x"5351", 
    x"534e", x"534c", x"534a", x"5347", x"5345", x"5342", x"5340", x"533e", 
    x"533b", x"5339", x"5336", x"5334", x"5332", x"532f", x"532d", x"532a", 
    x"5328", x"5326", x"5323", x"5321", x"531f", x"531c", x"531a", x"5317", 
    x"5315", x"5313", x"5310", x"530e", x"530b", x"5309", x"5307", x"5304", 
    x"5302", x"52ff", x"52fd", x"52fb", x"52f8", x"52f6", x"52f4", x"52f1", 
    x"52ef", x"52ec", x"52ea", x"52e8", x"52e5", x"52e3", x"52e0", x"52de", 
    x"52dc", x"52d9", x"52d7", x"52d4", x"52d2", x"52d0", x"52cd", x"52cb", 
    x"52c8", x"52c6", x"52c4", x"52c1", x"52bf", x"52bc", x"52ba", x"52b8", 
    x"52b5", x"52b3", x"52b0", x"52ae", x"52ac", x"52a9", x"52a7", x"52a4", 
    x"52a2", x"52a0", x"529d", x"529b", x"5298", x"5296", x"5294", x"5291", 
    x"528f", x"528c", x"528a", x"5288", x"5285", x"5283", x"5280", x"527e", 
    x"527c", x"5279", x"5277", x"5274", x"5272", x"5270", x"526d", x"526b", 
    x"5268", x"5266", x"5264", x"5261", x"525f", x"525c", x"525a", x"5258", 
    x"5255", x"5253", x"5250", x"524e", x"524c", x"5249", x"5247", x"5244", 
    x"5242", x"5240", x"523d", x"523b", x"5238", x"5236", x"5233", x"5231", 
    x"522f", x"522c", x"522a", x"5227", x"5225", x"5223", x"5220", x"521e", 
    x"521b", x"5219", x"5217", x"5214", x"5212", x"520f", x"520d", x"520b", 
    x"5208", x"5206", x"5203", x"5201", x"51fe", x"51fc", x"51fa", x"51f7", 
    x"51f5", x"51f2", x"51f0", x"51ee", x"51eb", x"51e9", x"51e6", x"51e4", 
    x"51e2", x"51df", x"51dd", x"51da", x"51d8", x"51d5", x"51d3", x"51d1", 
    x"51ce", x"51cc", x"51c9", x"51c7", x"51c5", x"51c2", x"51c0", x"51bd", 
    x"51bb", x"51b8", x"51b6", x"51b4", x"51b1", x"51af", x"51ac", x"51aa", 
    x"51a8", x"51a5", x"51a3", x"51a0", x"519e", x"519b", x"5199", x"5197", 
    x"5194", x"5192", x"518f", x"518d", x"518a", x"5188", x"5186", x"5183", 
    x"5181", x"517e", x"517c", x"517a", x"5177", x"5175", x"5172", x"5170", 
    x"516d", x"516b", x"5169", x"5166", x"5164", x"5161", x"515f", x"515c", 
    x"515a", x"5158", x"5155", x"5153", x"5150", x"514e", x"514b", x"5149", 
    x"5147", x"5144", x"5142", x"513f", x"513d", x"513a", x"5138", x"5136", 
    x"5133", x"5131", x"512e", x"512c", x"5129", x"5127", x"5125", x"5122", 
    x"5120", x"511d", x"511b", x"5118", x"5116", x"5114", x"5111", x"510f", 
    x"510c", x"510a", x"5107", x"5105", x"5103", x"5100", x"50fe", x"50fb", 
    x"50f9", x"50f6", x"50f4", x"50f2", x"50ef", x"50ed", x"50ea", x"50e8", 
    x"50e5", x"50e3", x"50e0", x"50de", x"50dc", x"50d9", x"50d7", x"50d4", 
    x"50d2", x"50cf", x"50cd", x"50cb", x"50c8", x"50c6", x"50c3", x"50c1", 
    x"50be", x"50bc", x"50ba", x"50b7", x"50b5", x"50b2", x"50b0", x"50ad", 
    x"50ab", x"50a8", x"50a6", x"50a4", x"50a1", x"509f", x"509c", x"509a", 
    x"5097", x"5095", x"5092", x"5090", x"508e", x"508b", x"5089", x"5086", 
    x"5084", x"5081", x"507f", x"507c", x"507a", x"5078", x"5075", x"5073", 
    x"5070", x"506e", x"506b", x"5069", x"5067", x"5064", x"5062", x"505f", 
    x"505d", x"505a", x"5058", x"5055", x"5053", x"5050", x"504e", x"504c", 
    x"5049", x"5047", x"5044", x"5042", x"503f", x"503d", x"503a", x"5038", 
    x"5036", x"5033", x"5031", x"502e", x"502c", x"5029", x"5027", x"5024", 
    x"5022", x"5020", x"501d", x"501b", x"5018", x"5016", x"5013", x"5011", 
    x"500e", x"500c", x"5009", x"5007", x"5005", x"5002", x"5000", x"4ffd", 
    x"4ffb", x"4ff8", x"4ff6", x"4ff3", x"4ff1", x"4fef", x"4fec", x"4fea", 
    x"4fe7", x"4fe5", x"4fe2", x"4fe0", x"4fdd", x"4fdb", x"4fd8", x"4fd6", 
    x"4fd4", x"4fd1", x"4fcf", x"4fcc", x"4fca", x"4fc7", x"4fc5", x"4fc2", 
    x"4fc0", x"4fbd", x"4fbb", x"4fb8", x"4fb6", x"4fb4", x"4fb1", x"4faf", 
    x"4fac", x"4faa", x"4fa7", x"4fa5", x"4fa2", x"4fa0", x"4f9d", x"4f9b", 
    x"4f99", x"4f96", x"4f94", x"4f91", x"4f8f", x"4f8c", x"4f8a", x"4f87", 
    x"4f85", x"4f82", x"4f80", x"4f7d", x"4f7b", x"4f79", x"4f76", x"4f74", 
    x"4f71", x"4f6f", x"4f6c", x"4f6a", x"4f67", x"4f65", x"4f62", x"4f60", 
    x"4f5d", x"4f5b", x"4f58", x"4f56", x"4f54", x"4f51", x"4f4f", x"4f4c", 
    x"4f4a", x"4f47", x"4f45", x"4f42", x"4f40", x"4f3d", x"4f3b", x"4f38", 
    x"4f36", x"4f33", x"4f31", x"4f2f", x"4f2c", x"4f2a", x"4f27", x"4f25", 
    x"4f22", x"4f20", x"4f1d", x"4f1b", x"4f18", x"4f16", x"4f13", x"4f11", 
    x"4f0e", x"4f0c", x"4f0a", x"4f07", x"4f05", x"4f02", x"4f00", x"4efd", 
    x"4efb", x"4ef8", x"4ef6", x"4ef3", x"4ef1", x"4eee", x"4eec", x"4ee9", 
    x"4ee7", x"4ee4", x"4ee2", x"4edf", x"4edd", x"4edb", x"4ed8", x"4ed6", 
    x"4ed3", x"4ed1", x"4ece", x"4ecc", x"4ec9", x"4ec7", x"4ec4", x"4ec2", 
    x"4ebf", x"4ebd", x"4eba", x"4eb8", x"4eb5", x"4eb3", x"4eb0", x"4eae", 
    x"4eab", x"4ea9", x"4ea7", x"4ea4", x"4ea2", x"4e9f", x"4e9d", x"4e9a", 
    x"4e98", x"4e95", x"4e93", x"4e90", x"4e8e", x"4e8b", x"4e89", x"4e86", 
    x"4e84", x"4e81", x"4e7f", x"4e7c", x"4e7a", x"4e77", x"4e75", x"4e72", 
    x"4e70", x"4e6d", x"4e6b", x"4e68", x"4e66", x"4e64", x"4e61", x"4e5f", 
    x"4e5c", x"4e5a", x"4e57", x"4e55", x"4e52", x"4e50", x"4e4d", x"4e4b", 
    x"4e48", x"4e46", x"4e43", x"4e41", x"4e3e", x"4e3c", x"4e39", x"4e37", 
    x"4e34", x"4e32", x"4e2f", x"4e2d", x"4e2a", x"4e28", x"4e25", x"4e23", 
    x"4e20", x"4e1e", x"4e1b", x"4e19", x"4e16", x"4e14", x"4e11", x"4e0f", 
    x"4e0d", x"4e0a", x"4e08", x"4e05", x"4e03", x"4e00", x"4dfe", x"4dfb", 
    x"4df9", x"4df6", x"4df4", x"4df1", x"4def", x"4dec", x"4dea", x"4de7", 
    x"4de5", x"4de2", x"4de0", x"4ddd", x"4ddb", x"4dd8", x"4dd6", x"4dd3", 
    x"4dd1", x"4dce", x"4dcc", x"4dc9", x"4dc7", x"4dc4", x"4dc2", x"4dbf", 
    x"4dbd", x"4dba", x"4db8", x"4db5", x"4db3", x"4db0", x"4dae", x"4dab", 
    x"4da9", x"4da6", x"4da4", x"4da1", x"4d9f", x"4d9c", x"4d9a", x"4d97", 
    x"4d95", x"4d92", x"4d90", x"4d8d", x"4d8b", x"4d88", x"4d86", x"4d83", 
    x"4d81", x"4d7e", x"4d7c", x"4d79", x"4d77", x"4d74", x"4d72", x"4d6f", 
    x"4d6d", x"4d6a", x"4d68", x"4d65", x"4d63", x"4d60", x"4d5e", x"4d5b", 
    x"4d59", x"4d56", x"4d54", x"4d51", x"4d4f", x"4d4c", x"4d4a", x"4d47", 
    x"4d45", x"4d42", x"4d40", x"4d3d", x"4d3b", x"4d38", x"4d36", x"4d33", 
    x"4d31", x"4d2e", x"4d2c", x"4d29", x"4d27", x"4d24", x"4d22", x"4d1f", 
    x"4d1d", x"4d1a", x"4d18", x"4d15", x"4d13", x"4d10", x"4d0e", x"4d0b", 
    x"4d09", x"4d06", x"4d04", x"4d01", x"4cff", x"4cfc", x"4cfa", x"4cf7", 
    x"4cf4", x"4cf2", x"4cef", x"4ced", x"4cea", x"4ce8", x"4ce5", x"4ce3", 
    x"4ce0", x"4cde", x"4cdb", x"4cd9", x"4cd6", x"4cd4", x"4cd1", x"4ccf", 
    x"4ccc", x"4cca", x"4cc7", x"4cc5", x"4cc2", x"4cc0", x"4cbd", x"4cbb", 
    x"4cb8", x"4cb6", x"4cb3", x"4cb1", x"4cae", x"4cac", x"4ca9", x"4ca7", 
    x"4ca4", x"4ca2", x"4c9f", x"4c9d", x"4c9a", x"4c97", x"4c95", x"4c92", 
    x"4c90", x"4c8d", x"4c8b", x"4c88", x"4c86", x"4c83", x"4c81", x"4c7e", 
    x"4c7c", x"4c79", x"4c77", x"4c74", x"4c72", x"4c6f", x"4c6d", x"4c6a", 
    x"4c68", x"4c65", x"4c63", x"4c60", x"4c5e", x"4c5b", x"4c59", x"4c56", 
    x"4c53", x"4c51", x"4c4e", x"4c4c", x"4c49", x"4c47", x"4c44", x"4c42", 
    x"4c3f", x"4c3d", x"4c3a", x"4c38", x"4c35", x"4c33", x"4c30", x"4c2e", 
    x"4c2b", x"4c29", x"4c26", x"4c24", x"4c21", x"4c1e", x"4c1c", x"4c19", 
    x"4c17", x"4c14", x"4c12", x"4c0f", x"4c0d", x"4c0a", x"4c08", x"4c05", 
    x"4c03", x"4c00", x"4bfe", x"4bfb", x"4bf9", x"4bf6", x"4bf4", x"4bf1", 
    x"4bee", x"4bec", x"4be9", x"4be7", x"4be4", x"4be2", x"4bdf", x"4bdd", 
    x"4bda", x"4bd8", x"4bd5", x"4bd3", x"4bd0", x"4bce", x"4bcb", x"4bc8", 
    x"4bc6", x"4bc3", x"4bc1", x"4bbe", x"4bbc", x"4bb9", x"4bb7", x"4bb4", 
    x"4bb2", x"4baf", x"4bad", x"4baa", x"4ba8", x"4ba5", x"4ba2", x"4ba0", 
    x"4b9d", x"4b9b", x"4b98", x"4b96", x"4b93", x"4b91", x"4b8e", x"4b8c", 
    x"4b89", x"4b87", x"4b84", x"4b82", x"4b7f", x"4b7c", x"4b7a", x"4b77", 
    x"4b75", x"4b72", x"4b70", x"4b6d", x"4b6b", x"4b68", x"4b66", x"4b63", 
    x"4b61", x"4b5e", x"4b5b", x"4b59", x"4b56", x"4b54", x"4b51", x"4b4f", 
    x"4b4c", x"4b4a", x"4b47", x"4b45", x"4b42", x"4b40", x"4b3d", x"4b3a", 
    x"4b38", x"4b35", x"4b33", x"4b30", x"4b2e", x"4b2b", x"4b29", x"4b26", 
    x"4b24", x"4b21", x"4b1e", x"4b1c", x"4b19", x"4b17", x"4b14", x"4b12", 
    x"4b0f", x"4b0d", x"4b0a", x"4b08", x"4b05", x"4b02", x"4b00", x"4afd", 
    x"4afb", x"4af8", x"4af6", x"4af3", x"4af1", x"4aee", x"4aec", x"4ae9", 
    x"4ae6", x"4ae4", x"4ae1", x"4adf", x"4adc", x"4ada", x"4ad7", x"4ad5", 
    x"4ad2", x"4ad0", x"4acd", x"4aca", x"4ac8", x"4ac5", x"4ac3", x"4ac0", 
    x"4abe", x"4abb", x"4ab9", x"4ab6", x"4ab3", x"4ab1", x"4aae", x"4aac", 
    x"4aa9", x"4aa7", x"4aa4", x"4aa2", x"4a9f", x"4a9d", x"4a9a", x"4a97", 
    x"4a95", x"4a92", x"4a90", x"4a8d", x"4a8b", x"4a88", x"4a86", x"4a83", 
    x"4a80", x"4a7e", x"4a7b", x"4a79", x"4a76", x"4a74", x"4a71", x"4a6f", 
    x"4a6c", x"4a69", x"4a67", x"4a64", x"4a62", x"4a5f", x"4a5d", x"4a5a", 
    x"4a58", x"4a55", x"4a52", x"4a50", x"4a4d", x"4a4b", x"4a48", x"4a46", 
    x"4a43", x"4a41", x"4a3e", x"4a3b", x"4a39", x"4a36", x"4a34", x"4a31", 
    x"4a2f", x"4a2c", x"4a29", x"4a27", x"4a24", x"4a22", x"4a1f", x"4a1d", 
    x"4a1a", x"4a18", x"4a15", x"4a12", x"4a10", x"4a0d", x"4a0b", x"4a08", 
    x"4a06", x"4a03", x"4a00", x"49fe", x"49fb", x"49f9", x"49f6", x"49f4", 
    x"49f1", x"49ef", x"49ec", x"49e9", x"49e7", x"49e4", x"49e2", x"49df", 
    x"49dd", x"49da", x"49d7", x"49d5", x"49d2", x"49d0", x"49cd", x"49cb", 
    x"49c8", x"49c5", x"49c3", x"49c0", x"49be", x"49bb", x"49b9", x"49b6", 
    x"49b4", x"49b1", x"49ae", x"49ac", x"49a9", x"49a7", x"49a4", x"49a2", 
    x"499f", x"499c", x"499a", x"4997", x"4995", x"4992", x"4990", x"498d", 
    x"498a", x"4988", x"4985", x"4983", x"4980", x"497e", x"497b", x"4978", 
    x"4976", x"4973", x"4971", x"496e", x"496c", x"4969", x"4966", x"4964", 
    x"4961", x"495f", x"495c", x"495a", x"4957", x"4954", x"4952", x"494f", 
    x"494d", x"494a", x"4947", x"4945", x"4942", x"4940", x"493d", x"493b", 
    x"4938", x"4935", x"4933", x"4930", x"492e", x"492b", x"4929", x"4926", 
    x"4923", x"4921", x"491e", x"491c", x"4919", x"4917", x"4914", x"4911", 
    x"490f", x"490c", x"490a", x"4907", x"4904", x"4902", x"48ff", x"48fd", 
    x"48fa", x"48f8", x"48f5", x"48f2", x"48f0", x"48ed", x"48eb", x"48e8", 
    x"48e5", x"48e3", x"48e0", x"48de", x"48db", x"48d9", x"48d6", x"48d3", 
    x"48d1", x"48ce", x"48cc", x"48c9", x"48c6", x"48c4", x"48c1", x"48bf", 
    x"48bc", x"48ba", x"48b7", x"48b4", x"48b2", x"48af", x"48ad", x"48aa", 
    x"48a7", x"48a5", x"48a2", x"48a0", x"489d", x"489b", x"4898", x"4895", 
    x"4893", x"4890", x"488e", x"488b", x"4888", x"4886", x"4883", x"4881", 
    x"487e", x"487b", x"4879", x"4876", x"4874", x"4871", x"486f", x"486c", 
    x"4869", x"4867", x"4864", x"4862", x"485f", x"485c", x"485a", x"4857", 
    x"4855", x"4852", x"484f", x"484d", x"484a", x"4848", x"4845", x"4842", 
    x"4840", x"483d", x"483b", x"4838", x"4835", x"4833", x"4830", x"482e", 
    x"482b", x"4829", x"4826", x"4823", x"4821", x"481e", x"481c", x"4819", 
    x"4816", x"4814", x"4811", x"480f", x"480c", x"4809", x"4807", x"4804", 
    x"4802", x"47ff", x"47fc", x"47fa", x"47f7", x"47f5", x"47f2", x"47ef", 
    x"47ed", x"47ea", x"47e8", x"47e5", x"47e2", x"47e0", x"47dd", x"47db", 
    x"47d8", x"47d5", x"47d3", x"47d0", x"47ce", x"47cb", x"47c8", x"47c6", 
    x"47c3", x"47c1", x"47be", x"47bb", x"47b9", x"47b6", x"47b4", x"47b1", 
    x"47ae", x"47ac", x"47a9", x"47a7", x"47a4", x"47a1", x"479f", x"479c", 
    x"479a", x"4797", x"4794", x"4792", x"478f", x"478d", x"478a", x"4787", 
    x"4785", x"4782", x"4780", x"477d", x"477a", x"4778", x"4775", x"4772", 
    x"4770", x"476d", x"476b", x"4768", x"4765", x"4763", x"4760", x"475e", 
    x"475b", x"4758", x"4756", x"4753", x"4751", x"474e", x"474b", x"4749", 
    x"4746", x"4744", x"4741", x"473e", x"473c", x"4739", x"4736", x"4734", 
    x"4731", x"472f", x"472c", x"4729", x"4727", x"4724", x"4722", x"471f", 
    x"471c", x"471a", x"4717", x"4715", x"4712", x"470f", x"470d", x"470a", 
    x"4707", x"4705", x"4702", x"4700", x"46fd", x"46fa", x"46f8", x"46f5", 
    x"46f3", x"46f0", x"46ed", x"46eb", x"46e8", x"46e5", x"46e3", x"46e0", 
    x"46de", x"46db", x"46d8", x"46d6", x"46d3", x"46d1", x"46ce", x"46cb", 
    x"46c9", x"46c6", x"46c3", x"46c1", x"46be", x"46bc", x"46b9", x"46b6", 
    x"46b4", x"46b1", x"46af", x"46ac", x"46a9", x"46a7", x"46a4", x"46a1", 
    x"469f", x"469c", x"469a", x"4697", x"4694", x"4692", x"468f", x"468c", 
    x"468a", x"4687", x"4685", x"4682", x"467f", x"467d", x"467a", x"4677", 
    x"4675", x"4672", x"4670", x"466d", x"466a", x"4668", x"4665", x"4662", 
    x"4660", x"465d", x"465b", x"4658", x"4655", x"4653", x"4650", x"464d", 
    x"464b", x"4648", x"4646", x"4643", x"4640", x"463e", x"463b", x"4638", 
    x"4636", x"4633", x"4631", x"462e", x"462b", x"4629", x"4626", x"4623", 
    x"4621", x"461e", x"461c", x"4619", x"4616", x"4614", x"4611", x"460e", 
    x"460c", x"4609", x"4607", x"4604", x"4601", x"45ff", x"45fc", x"45f9", 
    x"45f7", x"45f4", x"45f2", x"45ef", x"45ec", x"45ea", x"45e7", x"45e4", 
    x"45e2", x"45df", x"45dc", x"45da", x"45d7", x"45d5", x"45d2", x"45cf", 
    x"45cd", x"45ca", x"45c7", x"45c5", x"45c2", x"45bf", x"45bd", x"45ba", 
    x"45b8", x"45b5", x"45b2", x"45b0", x"45ad", x"45aa", x"45a8", x"45a5", 
    x"45a3", x"45a0", x"459d", x"459b", x"4598", x"4595", x"4593", x"4590", 
    x"458d", x"458b", x"4588", x"4586", x"4583", x"4580", x"457e", x"457b", 
    x"4578", x"4576", x"4573", x"4570", x"456e", x"456b", x"4568", x"4566", 
    x"4563", x"4561", x"455e", x"455b", x"4559", x"4556", x"4553", x"4551", 
    x"454e", x"454b", x"4549", x"4546", x"4544", x"4541", x"453e", x"453c", 
    x"4539", x"4536", x"4534", x"4531", x"452e", x"452c", x"4529", x"4526", 
    x"4524", x"4521", x"451f", x"451c", x"4519", x"4517", x"4514", x"4511", 
    x"450f", x"450c", x"4509", x"4507", x"4504", x"4501", x"44ff", x"44fc", 
    x"44f9", x"44f7", x"44f4", x"44f2", x"44ef", x"44ec", x"44ea", x"44e7", 
    x"44e4", x"44e2", x"44df", x"44dc", x"44da", x"44d7", x"44d4", x"44d2", 
    x"44cf", x"44cc", x"44ca", x"44c7", x"44c5", x"44c2", x"44bf", x"44bd", 
    x"44ba", x"44b7", x"44b5", x"44b2", x"44af", x"44ad", x"44aa", x"44a7", 
    x"44a5", x"44a2", x"449f", x"449d", x"449a", x"4497", x"4495", x"4492", 
    x"448f", x"448d", x"448a", x"4488", x"4485", x"4482", x"4480", x"447d", 
    x"447a", x"4478", x"4475", x"4472", x"4470", x"446d", x"446a", x"4468", 
    x"4465", x"4462", x"4460", x"445d", x"445a", x"4458", x"4455", x"4452", 
    x"4450", x"444d", x"444a", x"4448", x"4445", x"4442", x"4440", x"443d", 
    x"443b", x"4438", x"4435", x"4433", x"4430", x"442d", x"442b", x"4428", 
    x"4425", x"4423", x"4420", x"441d", x"441b", x"4418", x"4415", x"4413", 
    x"4410", x"440d", x"440b", x"4408", x"4405", x"4403", x"4400", x"43fd", 
    x"43fb", x"43f8", x"43f5", x"43f3", x"43f0", x"43ed", x"43eb", x"43e8", 
    x"43e5", x"43e3", x"43e0", x"43dd", x"43db", x"43d8", x"43d5", x"43d3", 
    x"43d0", x"43cd", x"43cb", x"43c8", x"43c5", x"43c3", x"43c0", x"43bd", 
    x"43bb", x"43b8", x"43b5", x"43b3", x"43b0", x"43ad", x"43ab", x"43a8", 
    x"43a5", x"43a3", x"43a0", x"439d", x"439b", x"4398", x"4395", x"4393", 
    x"4390", x"438d", x"438b", x"4388", x"4385", x"4383", x"4380", x"437d", 
    x"437b", x"4378", x"4375", x"4373", x"4370", x"436d", x"436b", x"4368", 
    x"4365", x"4363", x"4360", x"435d", x"435b", x"4358", x"4355", x"4353", 
    x"4350", x"434d", x"434b", x"4348", x"4345", x"4343", x"4340", x"433d", 
    x"433b", x"4338", x"4335", x"4333", x"4330", x"432d", x"432b", x"4328", 
    x"4325", x"4323", x"4320", x"431d", x"431b", x"4318", x"4315", x"4313", 
    x"4310", x"430d", x"430a", x"4308", x"4305", x"4302", x"4300", x"42fd", 
    x"42fa", x"42f8", x"42f5", x"42f2", x"42f0", x"42ed", x"42ea", x"42e8", 
    x"42e5", x"42e2", x"42e0", x"42dd", x"42da", x"42d8", x"42d5", x"42d2", 
    x"42d0", x"42cd", x"42ca", x"42c8", x"42c5", x"42c2", x"42bf", x"42bd", 
    x"42ba", x"42b7", x"42b5", x"42b2", x"42af", x"42ad", x"42aa", x"42a7", 
    x"42a5", x"42a2", x"429f", x"429d", x"429a", x"4297", x"4295", x"4292", 
    x"428f", x"428d", x"428a", x"4287", x"4284", x"4282", x"427f", x"427c", 
    x"427a", x"4277", x"4274", x"4272", x"426f", x"426c", x"426a", x"4267", 
    x"4264", x"4262", x"425f", x"425c", x"425a", x"4257", x"4254", x"4251", 
    x"424f", x"424c", x"4249", x"4247", x"4244", x"4241", x"423f", x"423c", 
    x"4239", x"4237", x"4234", x"4231", x"422f", x"422c", x"4229", x"4226", 
    x"4224", x"4221", x"421e", x"421c", x"4219", x"4216", x"4214", x"4211", 
    x"420e", x"420c", x"4209", x"4206", x"4203", x"4201", x"41fe", x"41fb", 
    x"41f9", x"41f6", x"41f3", x"41f1", x"41ee", x"41eb", x"41e9", x"41e6", 
    x"41e3", x"41e0", x"41de", x"41db", x"41d8", x"41d6", x"41d3", x"41d0", 
    x"41ce", x"41cb", x"41c8", x"41c6", x"41c3", x"41c0", x"41bd", x"41bb", 
    x"41b8", x"41b5", x"41b3", x"41b0", x"41ad", x"41ab", x"41a8", x"41a5", 
    x"41a2", x"41a0", x"419d", x"419a", x"4198", x"4195", x"4192", x"4190", 
    x"418d", x"418a", x"4187", x"4185", x"4182", x"417f", x"417d", x"417a", 
    x"4177", x"4175", x"4172", x"416f", x"416d", x"416a", x"4167", x"4164", 
    x"4162", x"415f", x"415c", x"415a", x"4157", x"4154", x"4151", x"414f", 
    x"414c", x"4149", x"4147", x"4144", x"4141", x"413f", x"413c", x"4139", 
    x"4136", x"4134", x"4131", x"412e", x"412c", x"4129", x"4126", x"4124", 
    x"4121", x"411e", x"411b", x"4119", x"4116", x"4113", x"4111", x"410e", 
    x"410b", x"4108", x"4106", x"4103", x"4100", x"40fe", x"40fb", x"40f8", 
    x"40f6", x"40f3", x"40f0", x"40ed", x"40eb", x"40e8", x"40e5", x"40e3", 
    x"40e0", x"40dd", x"40da", x"40d8", x"40d5", x"40d2", x"40d0", x"40cd", 
    x"40ca", x"40c8", x"40c5", x"40c2", x"40bf", x"40bd", x"40ba", x"40b7", 
    x"40b5", x"40b2", x"40af", x"40ac", x"40aa", x"40a7", x"40a4", x"40a2", 
    x"409f", x"409c", x"4099", x"4097", x"4094", x"4091", x"408f", x"408c", 
    x"4089", x"4086", x"4084", x"4081", x"407e", x"407c", x"4079", x"4076", 
    x"4073", x"4071", x"406e", x"406b", x"4069", x"4066", x"4063", x"4060", 
    x"405e", x"405b", x"4058", x"4056", x"4053", x"4050", x"404d", x"404b", 
    x"4048", x"4045", x"4043", x"4040", x"403d", x"403a", x"4038", x"4035", 
    x"4032", x"4030", x"402d", x"402a", x"4027", x"4025", x"4022", x"401f", 
    x"401d", x"401a", x"4017", x"4014", x"4012", x"400f", x"400c", x"4009", 
    x"4007", x"4004", x"4001", x"3fff", x"3ffc", x"3ff9", x"3ff6", x"3ff4", 
    x"3ff1", x"3fee", x"3fec", x"3fe9", x"3fe6", x"3fe3", x"3fe1", x"3fde", 
    x"3fdb", x"3fd8", x"3fd6", x"3fd3", x"3fd0", x"3fce", x"3fcb", x"3fc8", 
    x"3fc5", x"3fc3", x"3fc0", x"3fbd", x"3fbb", x"3fb8", x"3fb5", x"3fb2", 
    x"3fb0", x"3fad", x"3faa", x"3fa7", x"3fa5", x"3fa2", x"3f9f", x"3f9d", 
    x"3f9a", x"3f97", x"3f94", x"3f92", x"3f8f", x"3f8c", x"3f89", x"3f87", 
    x"3f84", x"3f81", x"3f7f", x"3f7c", x"3f79", x"3f76", x"3f74", x"3f71", 
    x"3f6e", x"3f6b", x"3f69", x"3f66", x"3f63", x"3f61", x"3f5e", x"3f5b", 
    x"3f58", x"3f56", x"3f53", x"3f50", x"3f4d", x"3f4b", x"3f48", x"3f45", 
    x"3f43", x"3f40", x"3f3d", x"3f3a", x"3f38", x"3f35", x"3f32", x"3f2f", 
    x"3f2d", x"3f2a", x"3f27", x"3f24", x"3f22", x"3f1f", x"3f1c", x"3f1a", 
    x"3f17", x"3f14", x"3f11", x"3f0f", x"3f0c", x"3f09", x"3f06", x"3f04", 
    x"3f01", x"3efe", x"3efb", x"3ef9", x"3ef6", x"3ef3", x"3ef1", x"3eee", 
    x"3eeb", x"3ee8", x"3ee6", x"3ee3", x"3ee0", x"3edd", x"3edb", x"3ed8", 
    x"3ed5", x"3ed2", x"3ed0", x"3ecd", x"3eca", x"3ec7", x"3ec5", x"3ec2", 
    x"3ebf", x"3ebd", x"3eba", x"3eb7", x"3eb4", x"3eb2", x"3eaf", x"3eac", 
    x"3ea9", x"3ea7", x"3ea4", x"3ea1", x"3e9e", x"3e9c", x"3e99", x"3e96", 
    x"3e93", x"3e91", x"3e8e", x"3e8b", x"3e88", x"3e86", x"3e83", x"3e80", 
    x"3e7d", x"3e7b", x"3e78", x"3e75", x"3e73", x"3e70", x"3e6d", x"3e6a", 
    x"3e68", x"3e65", x"3e62", x"3e5f", x"3e5d", x"3e5a", x"3e57", x"3e54", 
    x"3e52", x"3e4f", x"3e4c", x"3e49", x"3e47", x"3e44", x"3e41", x"3e3e", 
    x"3e3c", x"3e39", x"3e36", x"3e33", x"3e31", x"3e2e", x"3e2b", x"3e28", 
    x"3e26", x"3e23", x"3e20", x"3e1d", x"3e1b", x"3e18", x"3e15", x"3e12", 
    x"3e10", x"3e0d", x"3e0a", x"3e07", x"3e05", x"3e02", x"3dff", x"3dfc", 
    x"3dfa", x"3df7", x"3df4", x"3df1", x"3def", x"3dec", x"3de9", x"3de6", 
    x"3de4", x"3de1", x"3dde", x"3ddb", x"3dd9", x"3dd6", x"3dd3", x"3dd0", 
    x"3dce", x"3dcb", x"3dc8", x"3dc5", x"3dc3", x"3dc0", x"3dbd", x"3dba", 
    x"3db8", x"3db5", x"3db2", x"3daf", x"3dad", x"3daa", x"3da7", x"3da4", 
    x"3da2", x"3d9f", x"3d9c", x"3d99", x"3d97", x"3d94", x"3d91", x"3d8e", 
    x"3d8c", x"3d89", x"3d86", x"3d83", x"3d81", x"3d7e", x"3d7b", x"3d78", 
    x"3d76", x"3d73", x"3d70", x"3d6d", x"3d6b", x"3d68", x"3d65", x"3d62", 
    x"3d60", x"3d5d", x"3d5a", x"3d57", x"3d55", x"3d52", x"3d4f", x"3d4c", 
    x"3d4a", x"3d47", x"3d44", x"3d41", x"3d3e", x"3d3c", x"3d39", x"3d36", 
    x"3d33", x"3d31", x"3d2e", x"3d2b", x"3d28", x"3d26", x"3d23", x"3d20", 
    x"3d1d", x"3d1b", x"3d18", x"3d15", x"3d12", x"3d10", x"3d0d", x"3d0a", 
    x"3d07", x"3d05", x"3d02", x"3cff", x"3cfc", x"3cf9", x"3cf7", x"3cf4", 
    x"3cf1", x"3cee", x"3cec", x"3ce9", x"3ce6", x"3ce3", x"3ce1", x"3cde", 
    x"3cdb", x"3cd8", x"3cd6", x"3cd3", x"3cd0", x"3ccd", x"3cca", x"3cc8", 
    x"3cc5", x"3cc2", x"3cbf", x"3cbd", x"3cba", x"3cb7", x"3cb4", x"3cb2", 
    x"3caf", x"3cac", x"3ca9", x"3ca7", x"3ca4", x"3ca1", x"3c9e", x"3c9b", 
    x"3c99", x"3c96", x"3c93", x"3c90", x"3c8e", x"3c8b", x"3c88", x"3c85", 
    x"3c83", x"3c80", x"3c7d", x"3c7a", x"3c77", x"3c75", x"3c72", x"3c6f", 
    x"3c6c", x"3c6a", x"3c67", x"3c64", x"3c61", x"3c5f", x"3c5c", x"3c59", 
    x"3c56", x"3c53", x"3c51", x"3c4e", x"3c4b", x"3c48", x"3c46", x"3c43", 
    x"3c40", x"3c3d", x"3c3b", x"3c38", x"3c35", x"3c32", x"3c2f", x"3c2d", 
    x"3c2a", x"3c27", x"3c24", x"3c22", x"3c1f", x"3c1c", x"3c19", x"3c16", 
    x"3c14", x"3c11", x"3c0e", x"3c0b", x"3c09", x"3c06", x"3c03", x"3c00", 
    x"3bfe", x"3bfb", x"3bf8", x"3bf5", x"3bf2", x"3bf0", x"3bed", x"3bea", 
    x"3be7", x"3be5", x"3be2", x"3bdf", x"3bdc", x"3bd9", x"3bd7", x"3bd4", 
    x"3bd1", x"3bce", x"3bcc", x"3bc9", x"3bc6", x"3bc3", x"3bc0", x"3bbe", 
    x"3bbb", x"3bb8", x"3bb5", x"3bb3", x"3bb0", x"3bad", x"3baa", x"3ba7", 
    x"3ba5", x"3ba2", x"3b9f", x"3b9c", x"3b9a", x"3b97", x"3b94", x"3b91", 
    x"3b8e", x"3b8c", x"3b89", x"3b86", x"3b83", x"3b81", x"3b7e", x"3b7b", 
    x"3b78", x"3b75", x"3b73", x"3b70", x"3b6d", x"3b6a", x"3b67", x"3b65", 
    x"3b62", x"3b5f", x"3b5c", x"3b5a", x"3b57", x"3b54", x"3b51", x"3b4e", 
    x"3b4c", x"3b49", x"3b46", x"3b43", x"3b40", x"3b3e", x"3b3b", x"3b38", 
    x"3b35", x"3b33", x"3b30", x"3b2d", x"3b2a", x"3b27", x"3b25", x"3b22", 
    x"3b1f", x"3b1c", x"3b19", x"3b17", x"3b14", x"3b11", x"3b0e", x"3b0c", 
    x"3b09", x"3b06", x"3b03", x"3b00", x"3afe", x"3afb", x"3af8", x"3af5", 
    x"3af2", x"3af0", x"3aed", x"3aea", x"3ae7", x"3ae5", x"3ae2", x"3adf", 
    x"3adc", x"3ad9", x"3ad7", x"3ad4", x"3ad1", x"3ace", x"3acb", x"3ac9", 
    x"3ac6", x"3ac3", x"3ac0", x"3abd", x"3abb", x"3ab8", x"3ab5", x"3ab2", 
    x"3ab0", x"3aad", x"3aaa", x"3aa7", x"3aa4", x"3aa2", x"3a9f", x"3a9c", 
    x"3a99", x"3a96", x"3a94", x"3a91", x"3a8e", x"3a8b", x"3a88", x"3a86", 
    x"3a83", x"3a80", x"3a7d", x"3a7a", x"3a78", x"3a75", x"3a72", x"3a6f", 
    x"3a6c", x"3a6a", x"3a67", x"3a64", x"3a61", x"3a5e", x"3a5c", x"3a59", 
    x"3a56", x"3a53", x"3a51", x"3a4e", x"3a4b", x"3a48", x"3a45", x"3a43", 
    x"3a40", x"3a3d", x"3a3a", x"3a37", x"3a35", x"3a32", x"3a2f", x"3a2c", 
    x"3a29", x"3a27", x"3a24", x"3a21", x"3a1e", x"3a1b", x"3a19", x"3a16", 
    x"3a13", x"3a10", x"3a0d", x"3a0b", x"3a08", x"3a05", x"3a02", x"39ff", 
    x"39fd", x"39fa", x"39f7", x"39f4", x"39f1", x"39ef", x"39ec", x"39e9", 
    x"39e6", x"39e3", x"39e1", x"39de", x"39db", x"39d8", x"39d5", x"39d3", 
    x"39d0", x"39cd", x"39ca", x"39c7", x"39c5", x"39c2", x"39bf", x"39bc", 
    x"39b9", x"39b6", x"39b4", x"39b1", x"39ae", x"39ab", x"39a8", x"39a6", 
    x"39a3", x"39a0", x"399d", x"399a", x"3998", x"3995", x"3992", x"398f", 
    x"398c", x"398a", x"3987", x"3984", x"3981", x"397e", x"397c", x"3979", 
    x"3976", x"3973", x"3970", x"396e", x"396b", x"3968", x"3965", x"3962", 
    x"3960", x"395d", x"395a", x"3957", x"3954", x"3951", x"394f", x"394c", 
    x"3949", x"3946", x"3943", x"3941", x"393e", x"393b", x"3938", x"3935", 
    x"3933", x"3930", x"392d", x"392a", x"3927", x"3924", x"3922", x"391f", 
    x"391c", x"3919", x"3916", x"3914", x"3911", x"390e", x"390b", x"3908", 
    x"3906", x"3903", x"3900", x"38fd", x"38fa", x"38f8", x"38f5", x"38f2", 
    x"38ef", x"38ec", x"38e9", x"38e7", x"38e4", x"38e1", x"38de", x"38db", 
    x"38d9", x"38d6", x"38d3", x"38d0", x"38cd", x"38ca", x"38c8", x"38c5", 
    x"38c2", x"38bf", x"38bc", x"38ba", x"38b7", x"38b4", x"38b1", x"38ae", 
    x"38ab", x"38a9", x"38a6", x"38a3", x"38a0", x"389d", x"389b", x"3898", 
    x"3895", x"3892", x"388f", x"388d", x"388a", x"3887", x"3884", x"3881", 
    x"387e", x"387c", x"3879", x"3876", x"3873", x"3870", x"386d", x"386b", 
    x"3868", x"3865", x"3862", x"385f", x"385d", x"385a", x"3857", x"3854", 
    x"3851", x"384e", x"384c", x"3849", x"3846", x"3843", x"3840", x"383e", 
    x"383b", x"3838", x"3835", x"3832", x"382f", x"382d", x"382a", x"3827", 
    x"3824", x"3821", x"381e", x"381c", x"3819", x"3816", x"3813", x"3810", 
    x"380e", x"380b", x"3808", x"3805", x"3802", x"37ff", x"37fd", x"37fa", 
    x"37f7", x"37f4", x"37f1", x"37ee", x"37ec", x"37e9", x"37e6", x"37e3", 
    x"37e0", x"37de", x"37db", x"37d8", x"37d5", x"37d2", x"37cf", x"37cd", 
    x"37ca", x"37c7", x"37c4", x"37c1", x"37be", x"37bc", x"37b9", x"37b6", 
    x"37b3", x"37b0", x"37ad", x"37ab", x"37a8", x"37a5", x"37a2", x"379f", 
    x"379c", x"379a", x"3797", x"3794", x"3791", x"378e", x"378b", x"3789", 
    x"3786", x"3783", x"3780", x"377d", x"377b", x"3778", x"3775", x"3772", 
    x"376f", x"376c", x"376a", x"3767", x"3764", x"3761", x"375e", x"375b", 
    x"3759", x"3756", x"3753", x"3750", x"374d", x"374a", x"3748", x"3745", 
    x"3742", x"373f", x"373c", x"3739", x"3737", x"3734", x"3731", x"372e", 
    x"372b", x"3728", x"3726", x"3723", x"3720", x"371d", x"371a", x"3717", 
    x"3715", x"3712", x"370f", x"370c", x"3709", x"3706", x"3703", x"3701", 
    x"36fe", x"36fb", x"36f8", x"36f5", x"36f2", x"36f0", x"36ed", x"36ea", 
    x"36e7", x"36e4", x"36e1", x"36df", x"36dc", x"36d9", x"36d6", x"36d3", 
    x"36d0", x"36ce", x"36cb", x"36c8", x"36c5", x"36c2", x"36bf", x"36bd", 
    x"36ba", x"36b7", x"36b4", x"36b1", x"36ae", x"36ab", x"36a9", x"36a6", 
    x"36a3", x"36a0", x"369d", x"369a", x"3698", x"3695", x"3692", x"368f", 
    x"368c", x"3689", x"3687", x"3684", x"3681", x"367e", x"367b", x"3678", 
    x"3676", x"3673", x"3670", x"366d", x"366a", x"3667", x"3664", x"3662", 
    x"365f", x"365c", x"3659", x"3656", x"3653", x"3651", x"364e", x"364b", 
    x"3648", x"3645", x"3642", x"363f", x"363d", x"363a", x"3637", x"3634", 
    x"3631", x"362e", x"362c", x"3629", x"3626", x"3623", x"3620", x"361d", 
    x"361a", x"3618", x"3615", x"3612", x"360f", x"360c", x"3609", x"3607", 
    x"3604", x"3601", x"35fe", x"35fb", x"35f8", x"35f5", x"35f3", x"35f0", 
    x"35ed", x"35ea", x"35e7", x"35e4", x"35e1", x"35df", x"35dc", x"35d9", 
    x"35d6", x"35d3", x"35d0", x"35ce", x"35cb", x"35c8", x"35c5", x"35c2", 
    x"35bf", x"35bc", x"35ba", x"35b7", x"35b4", x"35b1", x"35ae", x"35ab", 
    x"35a8", x"35a6", x"35a3", x"35a0", x"359d", x"359a", x"3597", x"3595", 
    x"3592", x"358f", x"358c", x"3589", x"3586", x"3583", x"3581", x"357e", 
    x"357b", x"3578", x"3575", x"3572", x"356f", x"356d", x"356a", x"3567", 
    x"3564", x"3561", x"355e", x"355b", x"3559", x"3556", x"3553", x"3550", 
    x"354d", x"354a", x"3547", x"3545", x"3542", x"353f", x"353c", x"3539", 
    x"3536", x"3533", x"3531", x"352e", x"352b", x"3528", x"3525", x"3522", 
    x"351f", x"351d", x"351a", x"3517", x"3514", x"3511", x"350e", x"350b", 
    x"3509", x"3506", x"3503", x"3500", x"34fd", x"34fa", x"34f7", x"34f5", 
    x"34f2", x"34ef", x"34ec", x"34e9", x"34e6", x"34e3", x"34e1", x"34de", 
    x"34db", x"34d8", x"34d5", x"34d2", x"34cf", x"34cc", x"34ca", x"34c7", 
    x"34c4", x"34c1", x"34be", x"34bb", x"34b8", x"34b6", x"34b3", x"34b0", 
    x"34ad", x"34aa", x"34a7", x"34a4", x"34a2", x"349f", x"349c", x"3499", 
    x"3496", x"3493", x"3490", x"348e", x"348b", x"3488", x"3485", x"3482", 
    x"347f", x"347c", x"3479", x"3477", x"3474", x"3471", x"346e", x"346b", 
    x"3468", x"3465", x"3463", x"3460", x"345d", x"345a", x"3457", x"3454", 
    x"3451", x"344e", x"344c", x"3449", x"3446", x"3443", x"3440", x"343d", 
    x"343a", x"3438", x"3435", x"3432", x"342f", x"342c", x"3429", x"3426", 
    x"3423", x"3421", x"341e", x"341b", x"3418", x"3415", x"3412", x"340f", 
    x"340c", x"340a", x"3407", x"3404", x"3401", x"33fe", x"33fb", x"33f8", 
    x"33f6", x"33f3", x"33f0", x"33ed", x"33ea", x"33e7", x"33e4", x"33e1", 
    x"33df", x"33dc", x"33d9", x"33d6", x"33d3", x"33d0", x"33cd", x"33ca", 
    x"33c8", x"33c5", x"33c2", x"33bf", x"33bc", x"33b9", x"33b6", x"33b3", 
    x"33b1", x"33ae", x"33ab", x"33a8", x"33a5", x"33a2", x"339f", x"339c", 
    x"339a", x"3397", x"3394", x"3391", x"338e", x"338b", x"3388", x"3385", 
    x"3383", x"3380", x"337d", x"337a", x"3377", x"3374", x"3371", x"336e", 
    x"336c", x"3369", x"3366", x"3363", x"3360", x"335d", x"335a", x"3357", 
    x"3355", x"3352", x"334f", x"334c", x"3349", x"3346", x"3343", x"3340", 
    x"333e", x"333b", x"3338", x"3335", x"3332", x"332f", x"332c", x"3329", 
    x"3326", x"3324", x"3321", x"331e", x"331b", x"3318", x"3315", x"3312", 
    x"330f", x"330d", x"330a", x"3307", x"3304", x"3301", x"32fe", x"32fb", 
    x"32f8", x"32f6", x"32f3", x"32f0", x"32ed", x"32ea", x"32e7", x"32e4", 
    x"32e1", x"32de", x"32dc", x"32d9", x"32d6", x"32d3", x"32d0", x"32cd", 
    x"32ca", x"32c7", x"32c5", x"32c2", x"32bf", x"32bc", x"32b9", x"32b6", 
    x"32b3", x"32b0", x"32ad", x"32ab", x"32a8", x"32a5", x"32a2", x"329f", 
    x"329c", x"3299", x"3296", x"3293", x"3291", x"328e", x"328b", x"3288", 
    x"3285", x"3282", x"327f", x"327c", x"3279", x"3277", x"3274", x"3271", 
    x"326e", x"326b", x"3268", x"3265", x"3262", x"325f", x"325d", x"325a", 
    x"3257", x"3254", x"3251", x"324e", x"324b", x"3248", x"3246", x"3243", 
    x"3240", x"323d", x"323a", x"3237", x"3234", x"3231", x"322e", x"322b", 
    x"3229", x"3226", x"3223", x"3220", x"321d", x"321a", x"3217", x"3214", 
    x"3211", x"320f", x"320c", x"3209", x"3206", x"3203", x"3200", x"31fd", 
    x"31fa", x"31f7", x"31f5", x"31f2", x"31ef", x"31ec", x"31e9", x"31e6", 
    x"31e3", x"31e0", x"31dd", x"31db", x"31d8", x"31d5", x"31d2", x"31cf", 
    x"31cc", x"31c9", x"31c6", x"31c3", x"31c0", x"31be", x"31bb", x"31b8", 
    x"31b5", x"31b2", x"31af", x"31ac", x"31a9", x"31a6", x"31a4", x"31a1", 
    x"319e", x"319b", x"3198", x"3195", x"3192", x"318f", x"318c", x"3189", 
    x"3187", x"3184", x"3181", x"317e", x"317b", x"3178", x"3175", x"3172", 
    x"316f", x"316c", x"316a", x"3167", x"3164", x"3161", x"315e", x"315b", 
    x"3158", x"3155", x"3152", x"3150", x"314d", x"314a", x"3147", x"3144", 
    x"3141", x"313e", x"313b", x"3138", x"3135", x"3133", x"3130", x"312d", 
    x"312a", x"3127", x"3124", x"3121", x"311e", x"311b", x"3118", x"3116", 
    x"3113", x"3110", x"310d", x"310a", x"3107", x"3104", x"3101", x"30fe", 
    x"30fb", x"30f8", x"30f6", x"30f3", x"30f0", x"30ed", x"30ea", x"30e7", 
    x"30e4", x"30e1", x"30de", x"30db", x"30d9", x"30d6", x"30d3", x"30d0", 
    x"30cd", x"30ca", x"30c7", x"30c4", x"30c1", x"30be", x"30bc", x"30b9", 
    x"30b6", x"30b3", x"30b0", x"30ad", x"30aa", x"30a7", x"30a4", x"30a1", 
    x"309e", x"309c", x"3099", x"3096", x"3093", x"3090", x"308d", x"308a", 
    x"3087", x"3084", x"3081", x"307e", x"307c", x"3079", x"3076", x"3073", 
    x"3070", x"306d", x"306a", x"3067", x"3064", x"3061", x"305e", x"305c", 
    x"3059", x"3056", x"3053", x"3050", x"304d", x"304a", x"3047", x"3044", 
    x"3041", x"303e", x"303c", x"3039", x"3036", x"3033", x"3030", x"302d", 
    x"302a", x"3027", x"3024", x"3021", x"301e", x"301c", x"3019", x"3016", 
    x"3013", x"3010", x"300d", x"300a", x"3007", x"3004", x"3001", x"2ffe", 
    x"2ffc", x"2ff9", x"2ff6", x"2ff3", x"2ff0", x"2fed", x"2fea", x"2fe7", 
    x"2fe4", x"2fe1", x"2fde", x"2fdb", x"2fd9", x"2fd6", x"2fd3", x"2fd0", 
    x"2fcd", x"2fca", x"2fc7", x"2fc4", x"2fc1", x"2fbe", x"2fbb", x"2fb9", 
    x"2fb6", x"2fb3", x"2fb0", x"2fad", x"2faa", x"2fa7", x"2fa4", x"2fa1", 
    x"2f9e", x"2f9b", x"2f98", x"2f96", x"2f93", x"2f90", x"2f8d", x"2f8a", 
    x"2f87", x"2f84", x"2f81", x"2f7e", x"2f7b", x"2f78", x"2f75", x"2f73", 
    x"2f70", x"2f6d", x"2f6a", x"2f67", x"2f64", x"2f61", x"2f5e", x"2f5b", 
    x"2f58", x"2f55", x"2f52", x"2f50", x"2f4d", x"2f4a", x"2f47", x"2f44", 
    x"2f41", x"2f3e", x"2f3b", x"2f38", x"2f35", x"2f32", x"2f2f", x"2f2c", 
    x"2f2a", x"2f27", x"2f24", x"2f21", x"2f1e", x"2f1b", x"2f18", x"2f15", 
    x"2f12", x"2f0f", x"2f0c", x"2f09", x"2f06", x"2f04", x"2f01", x"2efe", 
    x"2efb", x"2ef8", x"2ef5", x"2ef2", x"2eef", x"2eec", x"2ee9", x"2ee6", 
    x"2ee3", x"2ee1", x"2ede", x"2edb", x"2ed8", x"2ed5", x"2ed2", x"2ecf", 
    x"2ecc", x"2ec9", x"2ec6", x"2ec3", x"2ec0", x"2ebd", x"2eba", x"2eb8", 
    x"2eb5", x"2eb2", x"2eaf", x"2eac", x"2ea9", x"2ea6", x"2ea3", x"2ea0", 
    x"2e9d", x"2e9a", x"2e97", x"2e94", x"2e92", x"2e8f", x"2e8c", x"2e89", 
    x"2e86", x"2e83", x"2e80", x"2e7d", x"2e7a", x"2e77", x"2e74", x"2e71", 
    x"2e6e", x"2e6b", x"2e69", x"2e66", x"2e63", x"2e60", x"2e5d", x"2e5a", 
    x"2e57", x"2e54", x"2e51", x"2e4e", x"2e4b", x"2e48", x"2e45", x"2e42", 
    x"2e40", x"2e3d", x"2e3a", x"2e37", x"2e34", x"2e31", x"2e2e", x"2e2b", 
    x"2e28", x"2e25", x"2e22", x"2e1f", x"2e1c", x"2e19", x"2e17", x"2e14", 
    x"2e11", x"2e0e", x"2e0b", x"2e08", x"2e05", x"2e02", x"2dff", x"2dfc", 
    x"2df9", x"2df6", x"2df3", x"2df0", x"2dee", x"2deb", x"2de8", x"2de5", 
    x"2de2", x"2ddf", x"2ddc", x"2dd9", x"2dd6", x"2dd3", x"2dd0", x"2dcd", 
    x"2dca", x"2dc7", x"2dc4", x"2dc2", x"2dbf", x"2dbc", x"2db9", x"2db6", 
    x"2db3", x"2db0", x"2dad", x"2daa", x"2da7", x"2da4", x"2da1", x"2d9e", 
    x"2d9b", x"2d98", x"2d95", x"2d93", x"2d90", x"2d8d", x"2d8a", x"2d87", 
    x"2d84", x"2d81", x"2d7e", x"2d7b", x"2d78", x"2d75", x"2d72", x"2d6f", 
    x"2d6c", x"2d69", x"2d67", x"2d64", x"2d61", x"2d5e", x"2d5b", x"2d58", 
    x"2d55", x"2d52", x"2d4f", x"2d4c", x"2d49", x"2d46", x"2d43", x"2d40", 
    x"2d3d", x"2d3a", x"2d37", x"2d35", x"2d32", x"2d2f", x"2d2c", x"2d29", 
    x"2d26", x"2d23", x"2d20", x"2d1d", x"2d1a", x"2d17", x"2d14", x"2d11", 
    x"2d0e", x"2d0b", x"2d08", x"2d06", x"2d03", x"2d00", x"2cfd", x"2cfa", 
    x"2cf7", x"2cf4", x"2cf1", x"2cee", x"2ceb", x"2ce8", x"2ce5", x"2ce2", 
    x"2cdf", x"2cdc", x"2cd9", x"2cd6", x"2cd4", x"2cd1", x"2cce", x"2ccb", 
    x"2cc8", x"2cc5", x"2cc2", x"2cbf", x"2cbc", x"2cb9", x"2cb6", x"2cb3", 
    x"2cb0", x"2cad", x"2caa", x"2ca7", x"2ca4", x"2ca1", x"2c9f", x"2c9c", 
    x"2c99", x"2c96", x"2c93", x"2c90", x"2c8d", x"2c8a", x"2c87", x"2c84", 
    x"2c81", x"2c7e", x"2c7b", x"2c78", x"2c75", x"2c72", x"2c6f", x"2c6c", 
    x"2c6a", x"2c67", x"2c64", x"2c61", x"2c5e", x"2c5b", x"2c58", x"2c55", 
    x"2c52", x"2c4f", x"2c4c", x"2c49", x"2c46", x"2c43", x"2c40", x"2c3d", 
    x"2c3a", x"2c37", x"2c34", x"2c32", x"2c2f", x"2c2c", x"2c29", x"2c26", 
    x"2c23", x"2c20", x"2c1d", x"2c1a", x"2c17", x"2c14", x"2c11", x"2c0e", 
    x"2c0b", x"2c08", x"2c05", x"2c02", x"2bff", x"2bfc", x"2bf9", x"2bf7", 
    x"2bf4", x"2bf1", x"2bee", x"2beb", x"2be8", x"2be5", x"2be2", x"2bdf", 
    x"2bdc", x"2bd9", x"2bd6", x"2bd3", x"2bd0", x"2bcd", x"2bca", x"2bc7", 
    x"2bc4", x"2bc1", x"2bbe", x"2bbb", x"2bb9", x"2bb6", x"2bb3", x"2bb0", 
    x"2bad", x"2baa", x"2ba7", x"2ba4", x"2ba1", x"2b9e", x"2b9b", x"2b98", 
    x"2b95", x"2b92", x"2b8f", x"2b8c", x"2b89", x"2b86", x"2b83", x"2b80", 
    x"2b7d", x"2b7b", x"2b78", x"2b75", x"2b72", x"2b6f", x"2b6c", x"2b69", 
    x"2b66", x"2b63", x"2b60", x"2b5d", x"2b5a", x"2b57", x"2b54", x"2b51", 
    x"2b4e", x"2b4b", x"2b48", x"2b45", x"2b42", x"2b3f", x"2b3c", x"2b39", 
    x"2b37", x"2b34", x"2b31", x"2b2e", x"2b2b", x"2b28", x"2b25", x"2b22", 
    x"2b1f", x"2b1c", x"2b19", x"2b16", x"2b13", x"2b10", x"2b0d", x"2b0a", 
    x"2b07", x"2b04", x"2b01", x"2afe", x"2afb", x"2af8", x"2af5", x"2af2", 
    x"2af0", x"2aed", x"2aea", x"2ae7", x"2ae4", x"2ae1", x"2ade", x"2adb", 
    x"2ad8", x"2ad5", x"2ad2", x"2acf", x"2acc", x"2ac9", x"2ac6", x"2ac3", 
    x"2ac0", x"2abd", x"2aba", x"2ab7", x"2ab4", x"2ab1", x"2aae", x"2aab", 
    x"2aa8", x"2aa6", x"2aa3", x"2aa0", x"2a9d", x"2a9a", x"2a97", x"2a94", 
    x"2a91", x"2a8e", x"2a8b", x"2a88", x"2a85", x"2a82", x"2a7f", x"2a7c", 
    x"2a79", x"2a76", x"2a73", x"2a70", x"2a6d", x"2a6a", x"2a67", x"2a64", 
    x"2a61", x"2a5e", x"2a5b", x"2a58", x"2a56", x"2a53", x"2a50", x"2a4d", 
    x"2a4a", x"2a47", x"2a44", x"2a41", x"2a3e", x"2a3b", x"2a38", x"2a35", 
    x"2a32", x"2a2f", x"2a2c", x"2a29", x"2a26", x"2a23", x"2a20", x"2a1d", 
    x"2a1a", x"2a17", x"2a14", x"2a11", x"2a0e", x"2a0b", x"2a08", x"2a05", 
    x"2a02", x"29ff", x"29fd", x"29fa", x"29f7", x"29f4", x"29f1", x"29ee", 
    x"29eb", x"29e8", x"29e5", x"29e2", x"29df", x"29dc", x"29d9", x"29d6", 
    x"29d3", x"29d0", x"29cd", x"29ca", x"29c7", x"29c4", x"29c1", x"29be", 
    x"29bb", x"29b8", x"29b5", x"29b2", x"29af", x"29ac", x"29a9", x"29a6", 
    x"29a3", x"29a0", x"299e", x"299b", x"2998", x"2995", x"2992", x"298f", 
    x"298c", x"2989", x"2986", x"2983", x"2980", x"297d", x"297a", x"2977", 
    x"2974", x"2971", x"296e", x"296b", x"2968", x"2965", x"2962", x"295f", 
    x"295c", x"2959", x"2956", x"2953", x"2950", x"294d", x"294a", x"2947", 
    x"2944", x"2941", x"293e", x"293b", x"2938", x"2935", x"2932", x"2930", 
    x"292d", x"292a", x"2927", x"2924", x"2921", x"291e", x"291b", x"2918", 
    x"2915", x"2912", x"290f", x"290c", x"2909", x"2906", x"2903", x"2900", 
    x"28fd", x"28fa", x"28f7", x"28f4", x"28f1", x"28ee", x"28eb", x"28e8", 
    x"28e5", x"28e2", x"28df", x"28dc", x"28d9", x"28d6", x"28d3", x"28d0", 
    x"28cd", x"28ca", x"28c7", x"28c4", x"28c1", x"28be", x"28bb", x"28b8", 
    x"28b5", x"28b3", x"28b0", x"28ad", x"28aa", x"28a7", x"28a4", x"28a1", 
    x"289e", x"289b", x"2898", x"2895", x"2892", x"288f", x"288c", x"2889", 
    x"2886", x"2883", x"2880", x"287d", x"287a", x"2877", x"2874", x"2871", 
    x"286e", x"286b", x"2868", x"2865", x"2862", x"285f", x"285c", x"2859", 
    x"2856", x"2853", x"2850", x"284d", x"284a", x"2847", x"2844", x"2841", 
    x"283e", x"283b", x"2838", x"2835", x"2832", x"282f", x"282c", x"2829", 
    x"2826", x"2823", x"2820", x"281d", x"281a", x"2817", x"2815", x"2812", 
    x"280f", x"280c", x"2809", x"2806", x"2803", x"2800", x"27fd", x"27fa", 
    x"27f7", x"27f4", x"27f1", x"27ee", x"27eb", x"27e8", x"27e5", x"27e2", 
    x"27df", x"27dc", x"27d9", x"27d6", x"27d3", x"27d0", x"27cd", x"27ca", 
    x"27c7", x"27c4", x"27c1", x"27be", x"27bb", x"27b8", x"27b5", x"27b2", 
    x"27af", x"27ac", x"27a9", x"27a6", x"27a3", x"27a0", x"279d", x"279a", 
    x"2797", x"2794", x"2791", x"278e", x"278b", x"2788", x"2785", x"2782", 
    x"277f", x"277c", x"2779", x"2776", x"2773", x"2770", x"276d", x"276a", 
    x"2767", x"2764", x"2761", x"275e", x"275b", x"2758", x"2755", x"2752", 
    x"274f", x"274c", x"2749", x"2746", x"2743", x"2740", x"273d", x"273a", 
    x"2737", x"2734", x"2731", x"272f", x"272c", x"2729", x"2726", x"2723", 
    x"2720", x"271d", x"271a", x"2717", x"2714", x"2711", x"270e", x"270b", 
    x"2708", x"2705", x"2702", x"26ff", x"26fc", x"26f9", x"26f6", x"26f3", 
    x"26f0", x"26ed", x"26ea", x"26e7", x"26e4", x"26e1", x"26de", x"26db", 
    x"26d8", x"26d5", x"26d2", x"26cf", x"26cc", x"26c9", x"26c6", x"26c3", 
    x"26c0", x"26bd", x"26ba", x"26b7", x"26b4", x"26b1", x"26ae", x"26ab", 
    x"26a8", x"26a5", x"26a2", x"269f", x"269c", x"2699", x"2696", x"2693", 
    x"2690", x"268d", x"268a", x"2687", x"2684", x"2681", x"267e", x"267b", 
    x"2678", x"2675", x"2672", x"266f", x"266c", x"2669", x"2666", x"2663", 
    x"2660", x"265d", x"265a", x"2657", x"2654", x"2651", x"264e", x"264b", 
    x"2648", x"2645", x"2642", x"263f", x"263c", x"2639", x"2636", x"2633", 
    x"2630", x"262d", x"262a", x"2627", x"2624", x"2621", x"261e", x"261b", 
    x"2618", x"2615", x"2612", x"260f", x"260c", x"2609", x"2606", x"2603", 
    x"2600", x"25fd", x"25fa", x"25f7", x"25f4", x"25f1", x"25ee", x"25eb", 
    x"25e8", x"25e5", x"25e2", x"25df", x"25dc", x"25d9", x"25d6", x"25d3", 
    x"25d0", x"25cd", x"25ca", x"25c7", x"25c4", x"25c1", x"25be", x"25bb", 
    x"25b8", x"25b5", x"25b2", x"25af", x"25ac", x"25a9", x"25a6", x"25a3", 
    x"25a0", x"259d", x"259a", x"2597", x"2594", x"2591", x"258e", x"258b", 
    x"2588", x"2585", x"2582", x"257f", x"257c", x"2579", x"2576", x"2573", 
    x"2570", x"256d", x"256a", x"2567", x"2564", x"2561", x"255e", x"255b", 
    x"2558", x"2555", x"2552", x"254f", x"254c", x"2549", x"2546", x"2543", 
    x"2540", x"253d", x"253a", x"2537", x"2534", x"2531", x"252e", x"252b", 
    x"2528", x"2525", x"2522", x"251f", x"251c", x"2519", x"2516", x"2513", 
    x"2510", x"250d", x"250a", x"2507", x"2504", x"2501", x"24fe", x"24fb", 
    x"24f8", x"24f5", x"24f2", x"24ef", x"24ec", x"24e9", x"24e6", x"24e3", 
    x"24e0", x"24dd", x"24da", x"24d7", x"24d4", x"24d1", x"24ce", x"24cb", 
    x"24c8", x"24c5", x"24c1", x"24be", x"24bb", x"24b8", x"24b5", x"24b2", 
    x"24af", x"24ac", x"24a9", x"24a6", x"24a3", x"24a0", x"249d", x"249a", 
    x"2497", x"2494", x"2491", x"248e", x"248b", x"2488", x"2485", x"2482", 
    x"247f", x"247c", x"2479", x"2476", x"2473", x"2470", x"246d", x"246a", 
    x"2467", x"2464", x"2461", x"245e", x"245b", x"2458", x"2455", x"2452", 
    x"244f", x"244c", x"2449", x"2446", x"2443", x"2440", x"243d", x"243a", 
    x"2437", x"2434", x"2431", x"242e", x"242b", x"2428", x"2425", x"2422", 
    x"241f", x"241c", x"2419", x"2416", x"2413", x"2410", x"240d", x"240a", 
    x"2407", x"2404", x"2401", x"23fe", x"23fb", x"23f8", x"23f5", x"23f2", 
    x"23ef", x"23ec", x"23e9", x"23e6", x"23e3", x"23e0", x"23dd", x"23da", 
    x"23d7", x"23d4", x"23d0", x"23cd", x"23ca", x"23c7", x"23c4", x"23c1", 
    x"23be", x"23bb", x"23b8", x"23b5", x"23b2", x"23af", x"23ac", x"23a9", 
    x"23a6", x"23a3", x"23a0", x"239d", x"239a", x"2397", x"2394", x"2391", 
    x"238e", x"238b", x"2388", x"2385", x"2382", x"237f", x"237c", x"2379", 
    x"2376", x"2373", x"2370", x"236d", x"236a", x"2367", x"2364", x"2361", 
    x"235e", x"235b", x"2358", x"2355", x"2352", x"234f", x"234c", x"2349", 
    x"2346", x"2343", x"2340", x"233d", x"233a", x"2337", x"2334", x"2331", 
    x"232e", x"232a", x"2327", x"2324", x"2321", x"231e", x"231b", x"2318", 
    x"2315", x"2312", x"230f", x"230c", x"2309", x"2306", x"2303", x"2300", 
    x"22fd", x"22fa", x"22f7", x"22f4", x"22f1", x"22ee", x"22eb", x"22e8", 
    x"22e5", x"22e2", x"22df", x"22dc", x"22d9", x"22d6", x"22d3", x"22d0", 
    x"22cd", x"22ca", x"22c7", x"22c4", x"22c1", x"22be", x"22bb", x"22b8", 
    x"22b5", x"22b2", x"22af", x"22ac", x"22a9", x"22a5", x"22a2", x"229f", 
    x"229c", x"2299", x"2296", x"2293", x"2290", x"228d", x"228a", x"2287", 
    x"2284", x"2281", x"227e", x"227b", x"2278", x"2275", x"2272", x"226f", 
    x"226c", x"2269", x"2266", x"2263", x"2260", x"225d", x"225a", x"2257", 
    x"2254", x"2251", x"224e", x"224b", x"2248", x"2245", x"2242", x"223f", 
    x"223c", x"2239", x"2236", x"2233", x"222f", x"222c", x"2229", x"2226", 
    x"2223", x"2220", x"221d", x"221a", x"2217", x"2214", x"2211", x"220e", 
    x"220b", x"2208", x"2205", x"2202", x"21ff", x"21fc", x"21f9", x"21f6", 
    x"21f3", x"21f0", x"21ed", x"21ea", x"21e7", x"21e4", x"21e1", x"21de", 
    x"21db", x"21d8", x"21d5", x"21d2", x"21cf", x"21cc", x"21c9", x"21c5", 
    x"21c2", x"21bf", x"21bc", x"21b9", x"21b6", x"21b3", x"21b0", x"21ad", 
    x"21aa", x"21a7", x"21a4", x"21a1", x"219e", x"219b", x"2198", x"2195", 
    x"2192", x"218f", x"218c", x"2189", x"2186", x"2183", x"2180", x"217d", 
    x"217a", x"2177", x"2174", x"2171", x"216e", x"216b", x"2168", x"2164", 
    x"2161", x"215e", x"215b", x"2158", x"2155", x"2152", x"214f", x"214c", 
    x"2149", x"2146", x"2143", x"2140", x"213d", x"213a", x"2137", x"2134", 
    x"2131", x"212e", x"212b", x"2128", x"2125", x"2122", x"211f", x"211c", 
    x"2119", x"2116", x"2113", x"2110", x"210c", x"2109", x"2106", x"2103", 
    x"2100", x"20fd", x"20fa", x"20f7", x"20f4", x"20f1", x"20ee", x"20eb", 
    x"20e8", x"20e5", x"20e2", x"20df", x"20dc", x"20d9", x"20d6", x"20d3", 
    x"20d0", x"20cd", x"20ca", x"20c7", x"20c4", x"20c1", x"20be", x"20bb", 
    x"20b7", x"20b4", x"20b1", x"20ae", x"20ab", x"20a8", x"20a5", x"20a2", 
    x"209f", x"209c", x"2099", x"2096", x"2093", x"2090", x"208d", x"208a", 
    x"2087", x"2084", x"2081", x"207e", x"207b", x"2078", x"2075", x"2072", 
    x"206f", x"206c", x"2068", x"2065", x"2062", x"205f", x"205c", x"2059", 
    x"2056", x"2053", x"2050", x"204d", x"204a", x"2047", x"2044", x"2041", 
    x"203e", x"203b", x"2038", x"2035", x"2032", x"202f", x"202c", x"2029", 
    x"2026", x"2023", x"2020", x"201c", x"2019", x"2016", x"2013", x"2010", 
    x"200d", x"200a", x"2007", x"2004", x"2001", x"1ffe", x"1ffb", x"1ff8", 
    x"1ff5", x"1ff2", x"1fef", x"1fec", x"1fe9", x"1fe6", x"1fe3", x"1fe0", 
    x"1fdd", x"1fda", x"1fd7", x"1fd3", x"1fd0", x"1fcd", x"1fca", x"1fc7", 
    x"1fc4", x"1fc1", x"1fbe", x"1fbb", x"1fb8", x"1fb5", x"1fb2", x"1faf", 
    x"1fac", x"1fa9", x"1fa6", x"1fa3", x"1fa0", x"1f9d", x"1f9a", x"1f97", 
    x"1f94", x"1f91", x"1f8d", x"1f8a", x"1f87", x"1f84", x"1f81", x"1f7e", 
    x"1f7b", x"1f78", x"1f75", x"1f72", x"1f6f", x"1f6c", x"1f69", x"1f66", 
    x"1f63", x"1f60", x"1f5d", x"1f5a", x"1f57", x"1f54", x"1f51", x"1f4e", 
    x"1f4a", x"1f47", x"1f44", x"1f41", x"1f3e", x"1f3b", x"1f38", x"1f35", 
    x"1f32", x"1f2f", x"1f2c", x"1f29", x"1f26", x"1f23", x"1f20", x"1f1d", 
    x"1f1a", x"1f17", x"1f14", x"1f11", x"1f0e", x"1f0a", x"1f07", x"1f04", 
    x"1f01", x"1efe", x"1efb", x"1ef8", x"1ef5", x"1ef2", x"1eef", x"1eec", 
    x"1ee9", x"1ee6", x"1ee3", x"1ee0", x"1edd", x"1eda", x"1ed7", x"1ed4", 
    x"1ed1", x"1ece", x"1eca", x"1ec7", x"1ec4", x"1ec1", x"1ebe", x"1ebb", 
    x"1eb8", x"1eb5", x"1eb2", x"1eaf", x"1eac", x"1ea9", x"1ea6", x"1ea3", 
    x"1ea0", x"1e9d", x"1e9a", x"1e97", x"1e94", x"1e91", x"1e8d", x"1e8a", 
    x"1e87", x"1e84", x"1e81", x"1e7e", x"1e7b", x"1e78", x"1e75", x"1e72", 
    x"1e6f", x"1e6c", x"1e69", x"1e66", x"1e63", x"1e60", x"1e5d", x"1e5a", 
    x"1e57", x"1e54", x"1e50", x"1e4d", x"1e4a", x"1e47", x"1e44", x"1e41", 
    x"1e3e", x"1e3b", x"1e38", x"1e35", x"1e32", x"1e2f", x"1e2c", x"1e29", 
    x"1e26", x"1e23", x"1e20", x"1e1d", x"1e19", x"1e16", x"1e13", x"1e10", 
    x"1e0d", x"1e0a", x"1e07", x"1e04", x"1e01", x"1dfe", x"1dfb", x"1df8", 
    x"1df5", x"1df2", x"1def", x"1dec", x"1de9", x"1de6", x"1de3", x"1ddf", 
    x"1ddc", x"1dd9", x"1dd6", x"1dd3", x"1dd0", x"1dcd", x"1dca", x"1dc7", 
    x"1dc4", x"1dc1", x"1dbe", x"1dbb", x"1db8", x"1db5", x"1db2", x"1daf", 
    x"1dac", x"1da8", x"1da5", x"1da2", x"1d9f", x"1d9c", x"1d99", x"1d96", 
    x"1d93", x"1d90", x"1d8d", x"1d8a", x"1d87", x"1d84", x"1d81", x"1d7e", 
    x"1d7b", x"1d78", x"1d75", x"1d71", x"1d6e", x"1d6b", x"1d68", x"1d65", 
    x"1d62", x"1d5f", x"1d5c", x"1d59", x"1d56", x"1d53", x"1d50", x"1d4d", 
    x"1d4a", x"1d47", x"1d44", x"1d41", x"1d3d", x"1d3a", x"1d37", x"1d34", 
    x"1d31", x"1d2e", x"1d2b", x"1d28", x"1d25", x"1d22", x"1d1f", x"1d1c", 
    x"1d19", x"1d16", x"1d13", x"1d10", x"1d0d", x"1d09", x"1d06", x"1d03", 
    x"1d00", x"1cfd", x"1cfa", x"1cf7", x"1cf4", x"1cf1", x"1cee", x"1ceb", 
    x"1ce8", x"1ce5", x"1ce2", x"1cdf", x"1cdc", x"1cd9", x"1cd5", x"1cd2", 
    x"1ccf", x"1ccc", x"1cc9", x"1cc6", x"1cc3", x"1cc0", x"1cbd", x"1cba", 
    x"1cb7", x"1cb4", x"1cb1", x"1cae", x"1cab", x"1ca8", x"1ca4", x"1ca1", 
    x"1c9e", x"1c9b", x"1c98", x"1c95", x"1c92", x"1c8f", x"1c8c", x"1c89", 
    x"1c86", x"1c83", x"1c80", x"1c7d", x"1c7a", x"1c77", x"1c73", x"1c70", 
    x"1c6d", x"1c6a", x"1c67", x"1c64", x"1c61", x"1c5e", x"1c5b", x"1c58", 
    x"1c55", x"1c52", x"1c4f", x"1c4c", x"1c49", x"1c46", x"1c42", x"1c3f", 
    x"1c3c", x"1c39", x"1c36", x"1c33", x"1c30", x"1c2d", x"1c2a", x"1c27", 
    x"1c24", x"1c21", x"1c1e", x"1c1b", x"1c18", x"1c14", x"1c11", x"1c0e", 
    x"1c0b", x"1c08", x"1c05", x"1c02", x"1bff", x"1bfc", x"1bf9", x"1bf6", 
    x"1bf3", x"1bf0", x"1bed", x"1bea", x"1be7", x"1be3", x"1be0", x"1bdd", 
    x"1bda", x"1bd7", x"1bd4", x"1bd1", x"1bce", x"1bcb", x"1bc8", x"1bc5", 
    x"1bc2", x"1bbf", x"1bbc", x"1bb9", x"1bb5", x"1bb2", x"1baf", x"1bac", 
    x"1ba9", x"1ba6", x"1ba3", x"1ba0", x"1b9d", x"1b9a", x"1b97", x"1b94", 
    x"1b91", x"1b8e", x"1b8a", x"1b87", x"1b84", x"1b81", x"1b7e", x"1b7b", 
    x"1b78", x"1b75", x"1b72", x"1b6f", x"1b6c", x"1b69", x"1b66", x"1b63", 
    x"1b60", x"1b5c", x"1b59", x"1b56", x"1b53", x"1b50", x"1b4d", x"1b4a", 
    x"1b47", x"1b44", x"1b41", x"1b3e", x"1b3b", x"1b38", x"1b35", x"1b31", 
    x"1b2e", x"1b2b", x"1b28", x"1b25", x"1b22", x"1b1f", x"1b1c", x"1b19", 
    x"1b16", x"1b13", x"1b10", x"1b0d", x"1b0a", x"1b07", x"1b03", x"1b00", 
    x"1afd", x"1afa", x"1af7", x"1af4", x"1af1", x"1aee", x"1aeb", x"1ae8", 
    x"1ae5", x"1ae2", x"1adf", x"1adc", x"1ad8", x"1ad5", x"1ad2", x"1acf", 
    x"1acc", x"1ac9", x"1ac6", x"1ac3", x"1ac0", x"1abd", x"1aba", x"1ab7", 
    x"1ab4", x"1ab1", x"1aad", x"1aaa", x"1aa7", x"1aa4", x"1aa1", x"1a9e", 
    x"1a9b", x"1a98", x"1a95", x"1a92", x"1a8f", x"1a8c", x"1a89", x"1a85", 
    x"1a82", x"1a7f", x"1a7c", x"1a79", x"1a76", x"1a73", x"1a70", x"1a6d", 
    x"1a6a", x"1a67", x"1a64", x"1a61", x"1a5e", x"1a5a", x"1a57", x"1a54", 
    x"1a51", x"1a4e", x"1a4b", x"1a48", x"1a45", x"1a42", x"1a3f", x"1a3c", 
    x"1a39", x"1a36", x"1a32", x"1a2f", x"1a2c", x"1a29", x"1a26", x"1a23", 
    x"1a20", x"1a1d", x"1a1a", x"1a17", x"1a14", x"1a11", x"1a0e", x"1a0b", 
    x"1a07", x"1a04", x"1a01", x"19fe", x"19fb", x"19f8", x"19f5", x"19f2", 
    x"19ef", x"19ec", x"19e9", x"19e6", x"19e3", x"19df", x"19dc", x"19d9", 
    x"19d6", x"19d3", x"19d0", x"19cd", x"19ca", x"19c7", x"19c4", x"19c1", 
    x"19be", x"19bb", x"19b7", x"19b4", x"19b1", x"19ae", x"19ab", x"19a8", 
    x"19a5", x"19a2", x"199f", x"199c", x"1999", x"1996", x"1993", x"198f", 
    x"198c", x"1989", x"1986", x"1983", x"1980", x"197d", x"197a", x"1977", 
    x"1974", x"1971", x"196e", x"196a", x"1967", x"1964", x"1961", x"195e", 
    x"195b", x"1958", x"1955", x"1952", x"194f", x"194c", x"1949", x"1946", 
    x"1942", x"193f", x"193c", x"1939", x"1936", x"1933", x"1930", x"192d", 
    x"192a", x"1927", x"1924", x"1921", x"191d", x"191a", x"1917", x"1914", 
    x"1911", x"190e", x"190b", x"1908", x"1905", x"1902", x"18ff", x"18fc", 
    x"18f9", x"18f5", x"18f2", x"18ef", x"18ec", x"18e9", x"18e6", x"18e3", 
    x"18e0", x"18dd", x"18da", x"18d7", x"18d4", x"18d0", x"18cd", x"18ca", 
    x"18c7", x"18c4", x"18c1", x"18be", x"18bb", x"18b8", x"18b5", x"18b2", 
    x"18af", x"18ab", x"18a8", x"18a5", x"18a2", x"189f", x"189c", x"1899", 
    x"1896", x"1893", x"1890", x"188d", x"188a", x"1886", x"1883", x"1880", 
    x"187d", x"187a", x"1877", x"1874", x"1871", x"186e", x"186b", x"1868", 
    x"1865", x"1861", x"185e", x"185b", x"1858", x"1855", x"1852", x"184f", 
    x"184c", x"1849", x"1846", x"1843", x"1840", x"183c", x"1839", x"1836", 
    x"1833", x"1830", x"182d", x"182a", x"1827", x"1824", x"1821", x"181e", 
    x"181b", x"1817", x"1814", x"1811", x"180e", x"180b", x"1808", x"1805", 
    x"1802", x"17ff", x"17fc", x"17f9", x"17f6", x"17f2", x"17ef", x"17ec", 
    x"17e9", x"17e6", x"17e3", x"17e0", x"17dd", x"17da", x"17d7", x"17d4", 
    x"17d0", x"17cd", x"17ca", x"17c7", x"17c4", x"17c1", x"17be", x"17bb", 
    x"17b8", x"17b5", x"17b2", x"17af", x"17ab", x"17a8", x"17a5", x"17a2", 
    x"179f", x"179c", x"1799", x"1796", x"1793", x"1790", x"178d", x"1789", 
    x"1786", x"1783", x"1780", x"177d", x"177a", x"1777", x"1774", x"1771", 
    x"176e", x"176b", x"1767", x"1764", x"1761", x"175e", x"175b", x"1758", 
    x"1755", x"1752", x"174f", x"174c", x"1749", x"1746", x"1742", x"173f", 
    x"173c", x"1739", x"1736", x"1733", x"1730", x"172d", x"172a", x"1727", 
    x"1724", x"1720", x"171d", x"171a", x"1717", x"1714", x"1711", x"170e", 
    x"170b", x"1708", x"1705", x"1702", x"16fe", x"16fb", x"16f8", x"16f5", 
    x"16f2", x"16ef", x"16ec", x"16e9", x"16e6", x"16e3", x"16e0", x"16dc", 
    x"16d9", x"16d6", x"16d3", x"16d0", x"16cd", x"16ca", x"16c7", x"16c4", 
    x"16c1", x"16be", x"16ba", x"16b7", x"16b4", x"16b1", x"16ae", x"16ab", 
    x"16a8", x"16a5", x"16a2", x"169f", x"169c", x"1698", x"1695", x"1692", 
    x"168f", x"168c", x"1689", x"1686", x"1683", x"1680", x"167d", x"167a", 
    x"1676", x"1673", x"1670", x"166d", x"166a", x"1667", x"1664", x"1661", 
    x"165e", x"165b", x"1657", x"1654", x"1651", x"164e", x"164b", x"1648", 
    x"1645", x"1642", x"163f", x"163c", x"1639", x"1635", x"1632", x"162f", 
    x"162c", x"1629", x"1626", x"1623", x"1620", x"161d", x"161a", x"1617", 
    x"1613", x"1610", x"160d", x"160a", x"1607", x"1604", x"1601", x"15fe", 
    x"15fb", x"15f8", x"15f4", x"15f1", x"15ee", x"15eb", x"15e8", x"15e5", 
    x"15e2", x"15df", x"15dc", x"15d9", x"15d6", x"15d2", x"15cf", x"15cc", 
    x"15c9", x"15c6", x"15c3", x"15c0", x"15bd", x"15ba", x"15b7", x"15b3", 
    x"15b0", x"15ad", x"15aa", x"15a7", x"15a4", x"15a1", x"159e", x"159b", 
    x"1598", x"1595", x"1591", x"158e", x"158b", x"1588", x"1585", x"1582", 
    x"157f", x"157c", x"1579", x"1576", x"1572", x"156f", x"156c", x"1569", 
    x"1566", x"1563", x"1560", x"155d", x"155a", x"1557", x"1553", x"1550", 
    x"154d", x"154a", x"1547", x"1544", x"1541", x"153e", x"153b", x"1538", 
    x"1534", x"1531", x"152e", x"152b", x"1528", x"1525", x"1522", x"151f", 
    x"151c", x"1519", x"1516", x"1512", x"150f", x"150c", x"1509", x"1506", 
    x"1503", x"1500", x"14fd", x"14fa", x"14f7", x"14f3", x"14f0", x"14ed", 
    x"14ea", x"14e7", x"14e4", x"14e1", x"14de", x"14db", x"14d8", x"14d4", 
    x"14d1", x"14ce", x"14cb", x"14c8", x"14c5", x"14c2", x"14bf", x"14bc", 
    x"14b9", x"14b5", x"14b2", x"14af", x"14ac", x"14a9", x"14a6", x"14a3", 
    x"14a0", x"149d", x"149a", x"1496", x"1493", x"1490", x"148d", x"148a", 
    x"1487", x"1484", x"1481", x"147e", x"147b", x"1477", x"1474", x"1471", 
    x"146e", x"146b", x"1468", x"1465", x"1462", x"145f", x"145c", x"1458", 
    x"1455", x"1452", x"144f", x"144c", x"1449", x"1446", x"1443", x"1440", 
    x"143c", x"1439", x"1436", x"1433", x"1430", x"142d", x"142a", x"1427", 
    x"1424", x"1421", x"141d", x"141a", x"1417", x"1414", x"1411", x"140e", 
    x"140b", x"1408", x"1405", x"1402", x"13fe", x"13fb", x"13f8", x"13f5", 
    x"13f2", x"13ef", x"13ec", x"13e9", x"13e6", x"13e3", x"13df", x"13dc", 
    x"13d9", x"13d6", x"13d3", x"13d0", x"13cd", x"13ca", x"13c7", x"13c3", 
    x"13c0", x"13bd", x"13ba", x"13b7", x"13b4", x"13b1", x"13ae", x"13ab", 
    x"13a8", x"13a4", x"13a1", x"139e", x"139b", x"1398", x"1395", x"1392", 
    x"138f", x"138c", x"1388", x"1385", x"1382", x"137f", x"137c", x"1379", 
    x"1376", x"1373", x"1370", x"136d", x"1369", x"1366", x"1363", x"1360", 
    x"135d", x"135a", x"1357", x"1354", x"1351", x"134d", x"134a", x"1347", 
    x"1344", x"1341", x"133e", x"133b", x"1338", x"1335", x"1332", x"132e", 
    x"132b", x"1328", x"1325", x"1322", x"131f", x"131c", x"1319", x"1316", 
    x"1312", x"130f", x"130c", x"1309", x"1306", x"1303", x"1300", x"12fd", 
    x"12fa", x"12f7", x"12f3", x"12f0", x"12ed", x"12ea", x"12e7", x"12e4", 
    x"12e1", x"12de", x"12db", x"12d7", x"12d4", x"12d1", x"12ce", x"12cb", 
    x"12c8", x"12c5", x"12c2", x"12bf", x"12bb", x"12b8", x"12b5", x"12b2", 
    x"12af", x"12ac", x"12a9", x"12a6", x"12a3", x"12a0", x"129c", x"1299", 
    x"1296", x"1293", x"1290", x"128d", x"128a", x"1287", x"1284", x"1280", 
    x"127d", x"127a", x"1277", x"1274", x"1271", x"126e", x"126b", x"1268", 
    x"1264", x"1261", x"125e", x"125b", x"1258", x"1255", x"1252", x"124f", 
    x"124c", x"1248", x"1245", x"1242", x"123f", x"123c", x"1239", x"1236", 
    x"1233", x"1230", x"122c", x"1229", x"1226", x"1223", x"1220", x"121d", 
    x"121a", x"1217", x"1214", x"1210", x"120d", x"120a", x"1207", x"1204", 
    x"1201", x"11fe", x"11fb", x"11f8", x"11f5", x"11f1", x"11ee", x"11eb", 
    x"11e8", x"11e5", x"11e2", x"11df", x"11dc", x"11d9", x"11d5", x"11d2", 
    x"11cf", x"11cc", x"11c9", x"11c6", x"11c3", x"11c0", x"11bd", x"11b9", 
    x"11b6", x"11b3", x"11b0", x"11ad", x"11aa", x"11a7", x"11a4", x"11a1", 
    x"119d", x"119a", x"1197", x"1194", x"1191", x"118e", x"118b", x"1188", 
    x"1185", x"1181", x"117e", x"117b", x"1178", x"1175", x"1172", x"116f", 
    x"116c", x"1168", x"1165", x"1162", x"115f", x"115c", x"1159", x"1156", 
    x"1153", x"1150", x"114c", x"1149", x"1146", x"1143", x"1140", x"113d", 
    x"113a", x"1137", x"1134", x"1130", x"112d", x"112a", x"1127", x"1124", 
    x"1121", x"111e", x"111b", x"1118", x"1114", x"1111", x"110e", x"110b", 
    x"1108", x"1105", x"1102", x"10ff", x"10fc", x"10f8", x"10f5", x"10f2", 
    x"10ef", x"10ec", x"10e9", x"10e6", x"10e3", x"10e0", x"10dc", x"10d9", 
    x"10d6", x"10d3", x"10d0", x"10cd", x"10ca", x"10c7", x"10c3", x"10c0", 
    x"10bd", x"10ba", x"10b7", x"10b4", x"10b1", x"10ae", x"10ab", x"10a7", 
    x"10a4", x"10a1", x"109e", x"109b", x"1098", x"1095", x"1092", x"108f", 
    x"108b", x"1088", x"1085", x"1082", x"107f", x"107c", x"1079", x"1076", 
    x"1072", x"106f", x"106c", x"1069", x"1066", x"1063", x"1060", x"105d", 
    x"105a", x"1056", x"1053", x"1050", x"104d", x"104a", x"1047", x"1044", 
    x"1041", x"103e", x"103a", x"1037", x"1034", x"1031", x"102e", x"102b", 
    x"1028", x"1025", x"1021", x"101e", x"101b", x"1018", x"1015", x"1012", 
    x"100f", x"100c", x"1009", x"1005", x"1002", x"0fff", x"0ffc", x"0ff9", 
    x"0ff6", x"0ff3", x"0ff0", x"0fec", x"0fe9", x"0fe6", x"0fe3", x"0fe0", 
    x"0fdd", x"0fda", x"0fd7", x"0fd4", x"0fd0", x"0fcd", x"0fca", x"0fc7", 
    x"0fc4", x"0fc1", x"0fbe", x"0fbb", x"0fb8", x"0fb4", x"0fb1", x"0fae", 
    x"0fab", x"0fa8", x"0fa5", x"0fa2", x"0f9f", x"0f9b", x"0f98", x"0f95", 
    x"0f92", x"0f8f", x"0f8c", x"0f89", x"0f86", x"0f82", x"0f7f", x"0f7c", 
    x"0f79", x"0f76", x"0f73", x"0f70", x"0f6d", x"0f6a", x"0f66", x"0f63", 
    x"0f60", x"0f5d", x"0f5a", x"0f57", x"0f54", x"0f51", x"0f4d", x"0f4a", 
    x"0f47", x"0f44", x"0f41", x"0f3e", x"0f3b", x"0f38", x"0f35", x"0f31", 
    x"0f2e", x"0f2b", x"0f28", x"0f25", x"0f22", x"0f1f", x"0f1c", x"0f18", 
    x"0f15", x"0f12", x"0f0f", x"0f0c", x"0f09", x"0f06", x"0f03", x"0eff", 
    x"0efc", x"0ef9", x"0ef6", x"0ef3", x"0ef0", x"0eed", x"0eea", x"0ee7", 
    x"0ee3", x"0ee0", x"0edd", x"0eda", x"0ed7", x"0ed4", x"0ed1", x"0ece", 
    x"0eca", x"0ec7", x"0ec4", x"0ec1", x"0ebe", x"0ebb", x"0eb8", x"0eb5", 
    x"0eb1", x"0eae", x"0eab", x"0ea8", x"0ea5", x"0ea2", x"0e9f", x"0e9c", 
    x"0e99", x"0e95", x"0e92", x"0e8f", x"0e8c", x"0e89", x"0e86", x"0e83", 
    x"0e80", x"0e7c", x"0e79", x"0e76", x"0e73", x"0e70", x"0e6d", x"0e6a", 
    x"0e67", x"0e63", x"0e60", x"0e5d", x"0e5a", x"0e57", x"0e54", x"0e51", 
    x"0e4e", x"0e4a", x"0e47", x"0e44", x"0e41", x"0e3e", x"0e3b", x"0e38", 
    x"0e35", x"0e32", x"0e2e", x"0e2b", x"0e28", x"0e25", x"0e22", x"0e1f", 
    x"0e1c", x"0e19", x"0e15", x"0e12", x"0e0f", x"0e0c", x"0e09", x"0e06", 
    x"0e03", x"0e00", x"0dfc", x"0df9", x"0df6", x"0df3", x"0df0", x"0ded", 
    x"0dea", x"0de7", x"0de3", x"0de0", x"0ddd", x"0dda", x"0dd7", x"0dd4", 
    x"0dd1", x"0dce", x"0dca", x"0dc7", x"0dc4", x"0dc1", x"0dbe", x"0dbb", 
    x"0db8", x"0db5", x"0db1", x"0dae", x"0dab", x"0da8", x"0da5", x"0da2", 
    x"0d9f", x"0d9c", x"0d98", x"0d95", x"0d92", x"0d8f", x"0d8c", x"0d89", 
    x"0d86", x"0d83", x"0d7f", x"0d7c", x"0d79", x"0d76", x"0d73", x"0d70", 
    x"0d6d", x"0d6a", x"0d66", x"0d63", x"0d60", x"0d5d", x"0d5a", x"0d57", 
    x"0d54", x"0d51", x"0d4e", x"0d4a", x"0d47", x"0d44", x"0d41", x"0d3e", 
    x"0d3b", x"0d38", x"0d35", x"0d31", x"0d2e", x"0d2b", x"0d28", x"0d25", 
    x"0d22", x"0d1f", x"0d1c", x"0d18", x"0d15", x"0d12", x"0d0f", x"0d0c", 
    x"0d09", x"0d06", x"0d03", x"0cff", x"0cfc", x"0cf9", x"0cf6", x"0cf3", 
    x"0cf0", x"0ced", x"0cea", x"0ce6", x"0ce3", x"0ce0", x"0cdd", x"0cda", 
    x"0cd7", x"0cd4", x"0cd1", x"0ccd", x"0cca", x"0cc7", x"0cc4", x"0cc1", 
    x"0cbe", x"0cbb", x"0cb7", x"0cb4", x"0cb1", x"0cae", x"0cab", x"0ca8", 
    x"0ca5", x"0ca2", x"0c9e", x"0c9b", x"0c98", x"0c95", x"0c92", x"0c8f", 
    x"0c8c", x"0c89", x"0c85", x"0c82", x"0c7f", x"0c7c", x"0c79", x"0c76", 
    x"0c73", x"0c70", x"0c6c", x"0c69", x"0c66", x"0c63", x"0c60", x"0c5d", 
    x"0c5a", x"0c57", x"0c53", x"0c50", x"0c4d", x"0c4a", x"0c47", x"0c44", 
    x"0c41", x"0c3e", x"0c3a", x"0c37", x"0c34", x"0c31", x"0c2e", x"0c2b", 
    x"0c28", x"0c25", x"0c21", x"0c1e", x"0c1b", x"0c18", x"0c15", x"0c12", 
    x"0c0f", x"0c0c", x"0c08", x"0c05", x"0c02", x"0bff", x"0bfc", x"0bf9", 
    x"0bf6", x"0bf3", x"0bef", x"0bec", x"0be9", x"0be6", x"0be3", x"0be0", 
    x"0bdd", x"0bd9", x"0bd6", x"0bd3", x"0bd0", x"0bcd", x"0bca", x"0bc7", 
    x"0bc4", x"0bc0", x"0bbd", x"0bba", x"0bb7", x"0bb4", x"0bb1", x"0bae", 
    x"0bab", x"0ba7", x"0ba4", x"0ba1", x"0b9e", x"0b9b", x"0b98", x"0b95", 
    x"0b92", x"0b8e", x"0b8b", x"0b88", x"0b85", x"0b82", x"0b7f", x"0b7c", 
    x"0b78", x"0b75", x"0b72", x"0b6f", x"0b6c", x"0b69", x"0b66", x"0b63", 
    x"0b5f", x"0b5c", x"0b59", x"0b56", x"0b53", x"0b50", x"0b4d", x"0b4a", 
    x"0b46", x"0b43", x"0b40", x"0b3d", x"0b3a", x"0b37", x"0b34", x"0b31", 
    x"0b2d", x"0b2a", x"0b27", x"0b24", x"0b21", x"0b1e", x"0b1b", x"0b17", 
    x"0b14", x"0b11", x"0b0e", x"0b0b", x"0b08", x"0b05", x"0b02", x"0afe", 
    x"0afb", x"0af8", x"0af5", x"0af2", x"0aef", x"0aec", x"0ae9", x"0ae5", 
    x"0ae2", x"0adf", x"0adc", x"0ad9", x"0ad6", x"0ad3", x"0acf", x"0acc", 
    x"0ac9", x"0ac6", x"0ac3", x"0ac0", x"0abd", x"0aba", x"0ab6", x"0ab3", 
    x"0ab0", x"0aad", x"0aaa", x"0aa7", x"0aa4", x"0aa1", x"0a9d", x"0a9a", 
    x"0a97", x"0a94", x"0a91", x"0a8e", x"0a8b", x"0a87", x"0a84", x"0a81", 
    x"0a7e", x"0a7b", x"0a78", x"0a75", x"0a72", x"0a6e", x"0a6b", x"0a68", 
    x"0a65", x"0a62", x"0a5f", x"0a5c", x"0a59", x"0a55", x"0a52", x"0a4f", 
    x"0a4c", x"0a49", x"0a46", x"0a43", x"0a3f", x"0a3c", x"0a39", x"0a36", 
    x"0a33", x"0a30", x"0a2d", x"0a2a", x"0a26", x"0a23", x"0a20", x"0a1d", 
    x"0a1a", x"0a17", x"0a14", x"0a11", x"0a0d", x"0a0a", x"0a07", x"0a04", 
    x"0a01", x"09fe", x"09fb", x"09f7", x"09f4", x"09f1", x"09ee", x"09eb", 
    x"09e8", x"09e5", x"09e2", x"09de", x"09db", x"09d8", x"09d5", x"09d2", 
    x"09cf", x"09cc", x"09c8", x"09c5", x"09c2", x"09bf", x"09bc", x"09b9", 
    x"09b6", x"09b3", x"09af", x"09ac", x"09a9", x"09a6", x"09a3", x"09a0", 
    x"099d", x"0999", x"0996", x"0993", x"0990", x"098d", x"098a", x"0987", 
    x"0984", x"0980", x"097d", x"097a", x"0977", x"0974", x"0971", x"096e", 
    x"096a", x"0967", x"0964", x"0961", x"095e", x"095b", x"0958", x"0955", 
    x"0951", x"094e", x"094b", x"0948", x"0945", x"0942", x"093f", x"093b", 
    x"0938", x"0935", x"0932", x"092f", x"092c", x"0929", x"0926", x"0922", 
    x"091f", x"091c", x"0919", x"0916", x"0913", x"0910", x"090c", x"0909", 
    x"0906", x"0903", x"0900", x"08fd", x"08fa", x"08f7", x"08f3", x"08f0", 
    x"08ed", x"08ea", x"08e7", x"08e4", x"08e1", x"08dd", x"08da", x"08d7", 
    x"08d4", x"08d1", x"08ce", x"08cb", x"08c8", x"08c4", x"08c1", x"08be", 
    x"08bb", x"08b8", x"08b5", x"08b2", x"08ae", x"08ab", x"08a8", x"08a5", 
    x"08a2", x"089f", x"089c", x"0899", x"0895", x"0892", x"088f", x"088c", 
    x"0889", x"0886", x"0883", x"087f", x"087c", x"0879", x"0876", x"0873", 
    x"0870", x"086d", x"086a", x"0866", x"0863", x"0860", x"085d", x"085a", 
    x"0857", x"0854", x"0850", x"084d", x"084a", x"0847", x"0844", x"0841", 
    x"083e", x"083a", x"0837", x"0834", x"0831", x"082e", x"082b", x"0828", 
    x"0825", x"0821", x"081e", x"081b", x"0818", x"0815", x"0812", x"080f", 
    x"080b", x"0808", x"0805", x"0802", x"07ff", x"07fc", x"07f9", x"07f6", 
    x"07f2", x"07ef", x"07ec", x"07e9", x"07e6", x"07e3", x"07e0", x"07dc", 
    x"07d9", x"07d6", x"07d3", x"07d0", x"07cd", x"07ca", x"07c6", x"07c3", 
    x"07c0", x"07bd", x"07ba", x"07b7", x"07b4", x"07b1", x"07ad", x"07aa", 
    x"07a7", x"07a4", x"07a1", x"079e", x"079b", x"0797", x"0794", x"0791", 
    x"078e", x"078b", x"0788", x"0785", x"0781", x"077e", x"077b", x"0778", 
    x"0775", x"0772", x"076f", x"076c", x"0768", x"0765", x"0762", x"075f", 
    x"075c", x"0759", x"0756", x"0752", x"074f", x"074c", x"0749", x"0746", 
    x"0743", x"0740", x"073c", x"0739", x"0736", x"0733", x"0730", x"072d", 
    x"072a", x"0727", x"0723", x"0720", x"071d", x"071a", x"0717", x"0714", 
    x"0711", x"070d", x"070a", x"0707", x"0704", x"0701", x"06fe", x"06fb", 
    x"06f7", x"06f4", x"06f1", x"06ee", x"06eb", x"06e8", x"06e5", x"06e2", 
    x"06de", x"06db", x"06d8", x"06d5", x"06d2", x"06cf", x"06cc", x"06c8", 
    x"06c5", x"06c2", x"06bf", x"06bc", x"06b9", x"06b6", x"06b2", x"06af", 
    x"06ac", x"06a9", x"06a6", x"06a3", x"06a0", x"069d", x"0699", x"0696", 
    x"0693", x"0690", x"068d", x"068a", x"0687", x"0683", x"0680", x"067d", 
    x"067a", x"0677", x"0674", x"0671", x"066d", x"066a", x"0667", x"0664", 
    x"0661", x"065e", x"065b", x"0657", x"0654", x"0651", x"064e", x"064b", 
    x"0648", x"0645", x"0642", x"063e", x"063b", x"0638", x"0635", x"0632", 
    x"062f", x"062c", x"0628", x"0625", x"0622", x"061f", x"061c", x"0619", 
    x"0616", x"0612", x"060f", x"060c", x"0609", x"0606", x"0603", x"0600", 
    x"05fc", x"05f9", x"05f6", x"05f3", x"05f0", x"05ed", x"05ea", x"05e7", 
    x"05e3", x"05e0", x"05dd", x"05da", x"05d7", x"05d4", x"05d1", x"05cd", 
    x"05ca", x"05c7", x"05c4", x"05c1", x"05be", x"05bb", x"05b7", x"05b4", 
    x"05b1", x"05ae", x"05ab", x"05a8", x"05a5", x"05a1", x"059e", x"059b", 
    x"0598", x"0595", x"0592", x"058f", x"058c", x"0588", x"0585", x"0582", 
    x"057f", x"057c", x"0579", x"0576", x"0572", x"056f", x"056c", x"0569", 
    x"0566", x"0563", x"0560", x"055c", x"0559", x"0556", x"0553", x"0550", 
    x"054d", x"054a", x"0546", x"0543", x"0540", x"053d", x"053a", x"0537", 
    x"0534", x"0530", x"052d", x"052a", x"0527", x"0524", x"0521", x"051e", 
    x"051b", x"0517", x"0514", x"0511", x"050e", x"050b", x"0508", x"0505", 
    x"0501", x"04fe", x"04fb", x"04f8", x"04f5", x"04f2", x"04ef", x"04eb", 
    x"04e8", x"04e5", x"04e2", x"04df", x"04dc", x"04d9", x"04d5", x"04d2", 
    x"04cf", x"04cc", x"04c9", x"04c6", x"04c3", x"04bf", x"04bc", x"04b9", 
    x"04b6", x"04b3", x"04b0", x"04ad", x"04aa", x"04a6", x"04a3", x"04a0", 
    x"049d", x"049a", x"0497", x"0494", x"0490", x"048d", x"048a", x"0487", 
    x"0484", x"0481", x"047e", x"047a", x"0477", x"0474", x"0471", x"046e", 
    x"046b", x"0468", x"0464", x"0461", x"045e", x"045b", x"0458", x"0455", 
    x"0452", x"044e", x"044b", x"0448", x"0445", x"0442", x"043f", x"043c", 
    x"0438", x"0435", x"0432", x"042f", x"042c", x"0429", x"0426", x"0423", 
    x"041f", x"041c", x"0419", x"0416", x"0413", x"0410", x"040d", x"0409", 
    x"0406", x"0403", x"0400", x"03fd", x"03fa", x"03f7", x"03f3", x"03f0", 
    x"03ed", x"03ea", x"03e7", x"03e4", x"03e1", x"03dd", x"03da", x"03d7", 
    x"03d4", x"03d1", x"03ce", x"03cb", x"03c7", x"03c4", x"03c1", x"03be", 
    x"03bb", x"03b8", x"03b5", x"03b1", x"03ae", x"03ab", x"03a8", x"03a5", 
    x"03a2", x"039f", x"039b", x"0398", x"0395", x"0392", x"038f", x"038c", 
    x"0389", x"0385", x"0382", x"037f", x"037c", x"0379", x"0376", x"0373", 
    x"0370", x"036c", x"0369", x"0366", x"0363", x"0360", x"035d", x"035a", 
    x"0356", x"0353", x"0350", x"034d", x"034a", x"0347", x"0344", x"0340", 
    x"033d", x"033a", x"0337", x"0334", x"0331", x"032e", x"032a", x"0327", 
    x"0324", x"0321", x"031e", x"031b", x"0318", x"0314", x"0311", x"030e", 
    x"030b", x"0308", x"0305", x"0302", x"02fe", x"02fb", x"02f8", x"02f5", 
    x"02f2", x"02ef", x"02ec", x"02e8", x"02e5", x"02e2", x"02df", x"02dc", 
    x"02d9", x"02d6", x"02d2", x"02cf", x"02cc", x"02c9", x"02c6", x"02c3", 
    x"02c0", x"02bd", x"02b9", x"02b6", x"02b3", x"02b0", x"02ad", x"02aa", 
    x"02a7", x"02a3", x"02a0", x"029d", x"029a", x"0297", x"0294", x"0291", 
    x"028d", x"028a", x"0287", x"0284", x"0281", x"027e", x"027b", x"0277", 
    x"0274", x"0271", x"026e", x"026b", x"0268", x"0265", x"0261", x"025e", 
    x"025b", x"0258", x"0255", x"0252", x"024f", x"024b", x"0248", x"0245", 
    x"0242", x"023f", x"023c", x"0239", x"0235", x"0232", x"022f", x"022c", 
    x"0229", x"0226", x"0223", x"021f", x"021c", x"0219", x"0216", x"0213", 
    x"0210", x"020d", x"0209", x"0206", x"0203", x"0200", x"01fd", x"01fa", 
    x"01f7", x"01f3", x"01f0", x"01ed", x"01ea", x"01e7", x"01e4", x"01e1", 
    x"01dd", x"01da", x"01d7", x"01d4", x"01d1", x"01ce", x"01cb", x"01c8", 
    x"01c4", x"01c1", x"01be", x"01bb", x"01b8", x"01b5", x"01b2", x"01ae", 
    x"01ab", x"01a8", x"01a5", x"01a2", x"019f", x"019c", x"0198", x"0195", 
    x"0192", x"018f", x"018c", x"0189", x"0186", x"0182", x"017f", x"017c", 
    x"0179", x"0176", x"0173", x"0170", x"016c", x"0169", x"0166", x"0163", 
    x"0160", x"015d", x"015a", x"0156", x"0153", x"0150", x"014d", x"014a", 
    x"0147", x"0144", x"0140", x"013d", x"013a", x"0137", x"0134", x"0131", 
    x"012e", x"012a", x"0127", x"0124", x"0121", x"011e", x"011b", x"0118", 
    x"0114", x"0111", x"010e", x"010b", x"0108", x"0105", x"0102", x"00fe", 
    x"00fb", x"00f8", x"00f5", x"00f2", x"00ef", x"00ec", x"00e8", x"00e5", 
    x"00e2", x"00df", x"00dc", x"00d9", x"00d6", x"00d2", x"00cf", x"00cc", 
    x"00c9", x"00c6", x"00c3", x"00c0", x"00bc", x"00b9", x"00b6", x"00b3", 
    x"00b0", x"00ad", x"00aa", x"00a6", x"00a3", x"00a0", x"009d", x"009a", 
    x"0097", x"0094", x"0091", x"008d", x"008a", x"0087", x"0084", x"0081", 
    x"007e", x"007b", x"0077", x"0074", x"0071", x"006e", x"006b", x"0068", 
    x"0065", x"0061", x"005e", x"005b", x"0058", x"0055", x"0052", x"004f", 
    x"004b", x"0048", x"0045", x"0042", x"003f", x"003c", x"0039", x"0035", 
    x"0032", x"002f", x"002c", x"0029", x"0026", x"0023", x"001f", x"001c", 
    x"0019", x"0016", x"0013", x"0010", x"000d", x"0009", x"0006", x"0003");

	constant icos : rom_mem :=( 
    x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", 
    x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", 
    x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", 
    x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", 
    x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", 
    x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", 
    x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", x"7fff", 
    x"7fff", x"7fff", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", 
    x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", 
    x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", 
    x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", 
    x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffe", 
    x"7ffe", x"7ffe", x"7ffe", x"7ffe", x"7ffd", x"7ffd", x"7ffd", x"7ffd", 
    x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", 
    x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", 
    x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", x"7ffd", 
    x"7ffd", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", 
    x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", 
    x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", x"7ffc", 
    x"7ffc", x"7ffb", x"7ffb", x"7ffb", x"7ffb", x"7ffb", x"7ffb", x"7ffb", 
    x"7ffb", x"7ffb", x"7ffb", x"7ffb", x"7ffb", x"7ffb", x"7ffb", x"7ffb", 
    x"7ffb", x"7ffb", x"7ffb", x"7ffb", x"7ffb", x"7ffa", x"7ffa", x"7ffa", 
    x"7ffa", x"7ffa", x"7ffa", x"7ffa", x"7ffa", x"7ffa", x"7ffa", x"7ffa", 
    x"7ffa", x"7ffa", x"7ffa", x"7ffa", x"7ffa", x"7ffa", x"7ffa", x"7ffa", 
    x"7ff9", x"7ff9", x"7ff9", x"7ff9", x"7ff9", x"7ff9", x"7ff9", x"7ff9", 
    x"7ff9", x"7ff9", x"7ff9", x"7ff9", x"7ff9", x"7ff9", x"7ff9", x"7ff9", 
    x"7ff8", x"7ff8", x"7ff8", x"7ff8", x"7ff8", x"7ff8", x"7ff8", x"7ff8", 
    x"7ff8", x"7ff8", x"7ff8", x"7ff8", x"7ff8", x"7ff8", x"7ff8", x"7ff8", 
    x"7ff7", x"7ff7", x"7ff7", x"7ff7", x"7ff7", x"7ff7", x"7ff7", x"7ff7", 
    x"7ff7", x"7ff7", x"7ff7", x"7ff7", x"7ff7", x"7ff7", x"7ff6", x"7ff6", 
    x"7ff6", x"7ff6", x"7ff6", x"7ff6", x"7ff6", x"7ff6", x"7ff6", x"7ff6", 
    x"7ff6", x"7ff6", x"7ff6", x"7ff6", x"7ff5", x"7ff5", x"7ff5", x"7ff5", 
    x"7ff5", x"7ff5", x"7ff5", x"7ff5", x"7ff5", x"7ff5", x"7ff5", x"7ff5", 
    x"7ff5", x"7ff4", x"7ff4", x"7ff4", x"7ff4", x"7ff4", x"7ff4", x"7ff4", 
    x"7ff4", x"7ff4", x"7ff4", x"7ff4", x"7ff4", x"7ff3", x"7ff3", x"7ff3", 
    x"7ff3", x"7ff3", x"7ff3", x"7ff3", x"7ff3", x"7ff3", x"7ff3", x"7ff3", 
    x"7ff3", x"7ff2", x"7ff2", x"7ff2", x"7ff2", x"7ff2", x"7ff2", x"7ff2", 
    x"7ff2", x"7ff2", x"7ff2", x"7ff2", x"7ff1", x"7ff1", x"7ff1", x"7ff1", 
    x"7ff1", x"7ff1", x"7ff1", x"7ff1", x"7ff1", x"7ff1", x"7ff1", x"7ff0", 
    x"7ff0", x"7ff0", x"7ff0", x"7ff0", x"7ff0", x"7ff0", x"7ff0", x"7ff0", 
    x"7ff0", x"7fef", x"7fef", x"7fef", x"7fef", x"7fef", x"7fef", x"7fef", 
    x"7fef", x"7fef", x"7fef", x"7fef", x"7fee", x"7fee", x"7fee", x"7fee", 
    x"7fee", x"7fee", x"7fee", x"7fee", x"7fee", x"7fed", x"7fed", x"7fed", 
    x"7fed", x"7fed", x"7fed", x"7fed", x"7fed", x"7fed", x"7fed", x"7fec", 
    x"7fec", x"7fec", x"7fec", x"7fec", x"7fec", x"7fec", x"7fec", x"7fec", 
    x"7feb", x"7feb", x"7feb", x"7feb", x"7feb", x"7feb", x"7feb", x"7feb", 
    x"7feb", x"7fea", x"7fea", x"7fea", x"7fea", x"7fea", x"7fea", x"7fea", 
    x"7fea", x"7fea", x"7fe9", x"7fe9", x"7fe9", x"7fe9", x"7fe9", x"7fe9", 
    x"7fe9", x"7fe9", x"7fe9", x"7fe8", x"7fe8", x"7fe8", x"7fe8", x"7fe8", 
    x"7fe8", x"7fe8", x"7fe8", x"7fe8", x"7fe7", x"7fe7", x"7fe7", x"7fe7", 
    x"7fe7", x"7fe7", x"7fe7", x"7fe7", x"7fe6", x"7fe6", x"7fe6", x"7fe6", 
    x"7fe6", x"7fe6", x"7fe6", x"7fe6", x"7fe5", x"7fe5", x"7fe5", x"7fe5", 
    x"7fe5", x"7fe5", x"7fe5", x"7fe5", x"7fe4", x"7fe4", x"7fe4", x"7fe4", 
    x"7fe4", x"7fe4", x"7fe4", x"7fe4", x"7fe3", x"7fe3", x"7fe3", x"7fe3", 
    x"7fe3", x"7fe3", x"7fe3", x"7fe3", x"7fe2", x"7fe2", x"7fe2", x"7fe2", 
    x"7fe2", x"7fe2", x"7fe2", x"7fe1", x"7fe1", x"7fe1", x"7fe1", x"7fe1", 
    x"7fe1", x"7fe1", x"7fe1", x"7fe0", x"7fe0", x"7fe0", x"7fe0", x"7fe0", 
    x"7fe0", x"7fe0", x"7fdf", x"7fdf", x"7fdf", x"7fdf", x"7fdf", x"7fdf", 
    x"7fdf", x"7fde", x"7fde", x"7fde", x"7fde", x"7fde", x"7fde", x"7fde", 
    x"7fdd", x"7fdd", x"7fdd", x"7fdd", x"7fdd", x"7fdd", x"7fdd", x"7fdc", 
    x"7fdc", x"7fdc", x"7fdc", x"7fdc", x"7fdc", x"7fdc", x"7fdb", x"7fdb", 
    x"7fdb", x"7fdb", x"7fdb", x"7fdb", x"7fdb", x"7fda", x"7fda", x"7fda", 
    x"7fda", x"7fda", x"7fda", x"7fda", x"7fd9", x"7fd9", x"7fd9", x"7fd9", 
    x"7fd9", x"7fd9", x"7fd8", x"7fd8", x"7fd8", x"7fd8", x"7fd8", x"7fd8", 
    x"7fd8", x"7fd7", x"7fd7", x"7fd7", x"7fd7", x"7fd7", x"7fd7", x"7fd6", 
    x"7fd6", x"7fd6", x"7fd6", x"7fd6", x"7fd6", x"7fd6", x"7fd5", x"7fd5", 
    x"7fd5", x"7fd5", x"7fd5", x"7fd5", x"7fd4", x"7fd4", x"7fd4", x"7fd4", 
    x"7fd4", x"7fd4", x"7fd3", x"7fd3", x"7fd3", x"7fd3", x"7fd3", x"7fd3", 
    x"7fd2", x"7fd2", x"7fd2", x"7fd2", x"7fd2", x"7fd2", x"7fd1", x"7fd1", 
    x"7fd1", x"7fd1", x"7fd1", x"7fd1", x"7fd0", x"7fd0", x"7fd0", x"7fd0", 
    x"7fd0", x"7fd0", x"7fcf", x"7fcf", x"7fcf", x"7fcf", x"7fcf", x"7fcf", 
    x"7fce", x"7fce", x"7fce", x"7fce", x"7fce", x"7fce", x"7fcd", x"7fcd", 
    x"7fcd", x"7fcd", x"7fcd", x"7fcd", x"7fcc", x"7fcc", x"7fcc", x"7fcc", 
    x"7fcc", x"7fcb", x"7fcb", x"7fcb", x"7fcb", x"7fcb", x"7fcb", x"7fca", 
    x"7fca", x"7fca", x"7fca", x"7fca", x"7fca", x"7fc9", x"7fc9", x"7fc9", 
    x"7fc9", x"7fc9", x"7fc8", x"7fc8", x"7fc8", x"7fc8", x"7fc8", x"7fc8", 
    x"7fc7", x"7fc7", x"7fc7", x"7fc7", x"7fc7", x"7fc6", x"7fc6", x"7fc6", 
    x"7fc6", x"7fc6", x"7fc6", x"7fc5", x"7fc5", x"7fc5", x"7fc5", x"7fc5", 
    x"7fc4", x"7fc4", x"7fc4", x"7fc4", x"7fc4", x"7fc3", x"7fc3", x"7fc3", 
    x"7fc3", x"7fc3", x"7fc2", x"7fc2", x"7fc2", x"7fc2", x"7fc2", x"7fc2", 
    x"7fc1", x"7fc1", x"7fc1", x"7fc1", x"7fc1", x"7fc0", x"7fc0", x"7fc0", 
    x"7fc0", x"7fc0", x"7fbf", x"7fbf", x"7fbf", x"7fbf", x"7fbf", x"7fbe", 
    x"7fbe", x"7fbe", x"7fbe", x"7fbe", x"7fbd", x"7fbd", x"7fbd", x"7fbd", 
    x"7fbd", x"7fbc", x"7fbc", x"7fbc", x"7fbc", x"7fbc", x"7fbb", x"7fbb", 
    x"7fbb", x"7fbb", x"7fbb", x"7fba", x"7fba", x"7fba", x"7fba", x"7fba", 
    x"7fb9", x"7fb9", x"7fb9", x"7fb9", x"7fb9", x"7fb8", x"7fb8", x"7fb8", 
    x"7fb8", x"7fb8", x"7fb7", x"7fb7", x"7fb7", x"7fb7", x"7fb6", x"7fb6", 
    x"7fb6", x"7fb6", x"7fb6", x"7fb5", x"7fb5", x"7fb5", x"7fb5", x"7fb5", 
    x"7fb4", x"7fb4", x"7fb4", x"7fb4", x"7fb4", x"7fb3", x"7fb3", x"7fb3", 
    x"7fb3", x"7fb2", x"7fb2", x"7fb2", x"7fb2", x"7fb2", x"7fb1", x"7fb1", 
    x"7fb1", x"7fb1", x"7fb1", x"7fb0", x"7fb0", x"7fb0", x"7fb0", x"7faf", 
    x"7faf", x"7faf", x"7faf", x"7faf", x"7fae", x"7fae", x"7fae", x"7fae", 
    x"7fad", x"7fad", x"7fad", x"7fad", x"7fad", x"7fac", x"7fac", x"7fac", 
    x"7fac", x"7fab", x"7fab", x"7fab", x"7fab", x"7fab", x"7faa", x"7faa", 
    x"7faa", x"7faa", x"7fa9", x"7fa9", x"7fa9", x"7fa9", x"7fa9", x"7fa8", 
    x"7fa8", x"7fa8", x"7fa8", x"7fa7", x"7fa7", x"7fa7", x"7fa7", x"7fa6", 
    x"7fa6", x"7fa6", x"7fa6", x"7fa6", x"7fa5", x"7fa5", x"7fa5", x"7fa5", 
    x"7fa4", x"7fa4", x"7fa4", x"7fa4", x"7fa3", x"7fa3", x"7fa3", x"7fa3", 
    x"7fa2", x"7fa2", x"7fa2", x"7fa2", x"7fa2", x"7fa1", x"7fa1", x"7fa1", 
    x"7fa1", x"7fa0", x"7fa0", x"7fa0", x"7fa0", x"7f9f", x"7f9f", x"7f9f", 
    x"7f9f", x"7f9e", x"7f9e", x"7f9e", x"7f9e", x"7f9d", x"7f9d", x"7f9d", 
    x"7f9d", x"7f9c", x"7f9c", x"7f9c", x"7f9c", x"7f9c", x"7f9b", x"7f9b", 
    x"7f9b", x"7f9b", x"7f9a", x"7f9a", x"7f9a", x"7f9a", x"7f99", x"7f99", 
    x"7f99", x"7f99", x"7f98", x"7f98", x"7f98", x"7f98", x"7f97", x"7f97", 
    x"7f97", x"7f97", x"7f96", x"7f96", x"7f96", x"7f96", x"7f95", x"7f95", 
    x"7f95", x"7f95", x"7f94", x"7f94", x"7f94", x"7f94", x"7f93", x"7f93", 
    x"7f93", x"7f93", x"7f92", x"7f92", x"7f92", x"7f91", x"7f91", x"7f91", 
    x"7f91", x"7f90", x"7f90", x"7f90", x"7f90", x"7f8f", x"7f8f", x"7f8f", 
    x"7f8f", x"7f8e", x"7f8e", x"7f8e", x"7f8e", x"7f8d", x"7f8d", x"7f8d", 
    x"7f8d", x"7f8c", x"7f8c", x"7f8c", x"7f8c", x"7f8b", x"7f8b", x"7f8b", 
    x"7f8a", x"7f8a", x"7f8a", x"7f8a", x"7f89", x"7f89", x"7f89", x"7f89", 
    x"7f88", x"7f88", x"7f88", x"7f88", x"7f87", x"7f87", x"7f87", x"7f86", 
    x"7f86", x"7f86", x"7f86", x"7f85", x"7f85", x"7f85", x"7f85", x"7f84", 
    x"7f84", x"7f84", x"7f83", x"7f83", x"7f83", x"7f83", x"7f82", x"7f82", 
    x"7f82", x"7f82", x"7f81", x"7f81", x"7f81", x"7f80", x"7f80", x"7f80", 
    x"7f80", x"7f7f", x"7f7f", x"7f7f", x"7f7f", x"7f7e", x"7f7e", x"7f7e", 
    x"7f7d", x"7f7d", x"7f7d", x"7f7d", x"7f7c", x"7f7c", x"7f7c", x"7f7b", 
    x"7f7b", x"7f7b", x"7f7b", x"7f7a", x"7f7a", x"7f7a", x"7f79", x"7f79", 
    x"7f79", x"7f79", x"7f78", x"7f78", x"7f78", x"7f77", x"7f77", x"7f77", 
    x"7f77", x"7f76", x"7f76", x"7f76", x"7f75", x"7f75", x"7f75", x"7f75", 
    x"7f74", x"7f74", x"7f74", x"7f73", x"7f73", x"7f73", x"7f73", x"7f72", 
    x"7f72", x"7f72", x"7f71", x"7f71", x"7f71", x"7f71", x"7f70", x"7f70", 
    x"7f70", x"7f6f", x"7f6f", x"7f6f", x"7f6e", x"7f6e", x"7f6e", x"7f6e", 
    x"7f6d", x"7f6d", x"7f6d", x"7f6c", x"7f6c", x"7f6c", x"7f6c", x"7f6b", 
    x"7f6b", x"7f6b", x"7f6a", x"7f6a", x"7f6a", x"7f69", x"7f69", x"7f69", 
    x"7f69", x"7f68", x"7f68", x"7f68", x"7f67", x"7f67", x"7f67", x"7f66", 
    x"7f66", x"7f66", x"7f65", x"7f65", x"7f65", x"7f65", x"7f64", x"7f64", 
    x"7f64", x"7f63", x"7f63", x"7f63", x"7f62", x"7f62", x"7f62", x"7f62", 
    x"7f61", x"7f61", x"7f61", x"7f60", x"7f60", x"7f60", x"7f5f", x"7f5f", 
    x"7f5f", x"7f5e", x"7f5e", x"7f5e", x"7f5e", x"7f5d", x"7f5d", x"7f5d", 
    x"7f5c", x"7f5c", x"7f5c", x"7f5b", x"7f5b", x"7f5b", x"7f5a", x"7f5a", 
    x"7f5a", x"7f59", x"7f59", x"7f59", x"7f58", x"7f58", x"7f58", x"7f58", 
    x"7f57", x"7f57", x"7f57", x"7f56", x"7f56", x"7f56", x"7f55", x"7f55", 
    x"7f55", x"7f54", x"7f54", x"7f54", x"7f53", x"7f53", x"7f53", x"7f52", 
    x"7f52", x"7f52", x"7f51", x"7f51", x"7f51", x"7f50", x"7f50", x"7f50", 
    x"7f50", x"7f4f", x"7f4f", x"7f4f", x"7f4e", x"7f4e", x"7f4e", x"7f4d", 
    x"7f4d", x"7f4d", x"7f4c", x"7f4c", x"7f4c", x"7f4b", x"7f4b", x"7f4b", 
    x"7f4a", x"7f4a", x"7f4a", x"7f49", x"7f49", x"7f49", x"7f48", x"7f48", 
    x"7f48", x"7f47", x"7f47", x"7f47", x"7f46", x"7f46", x"7f46", x"7f45", 
    x"7f45", x"7f45", x"7f44", x"7f44", x"7f44", x"7f43", x"7f43", x"7f43", 
    x"7f42", x"7f42", x"7f42", x"7f41", x"7f41", x"7f41", x"7f40", x"7f40", 
    x"7f40", x"7f3f", x"7f3f", x"7f3f", x"7f3e", x"7f3e", x"7f3e", x"7f3d", 
    x"7f3d", x"7f3d", x"7f3c", x"7f3c", x"7f3b", x"7f3b", x"7f3b", x"7f3a", 
    x"7f3a", x"7f3a", x"7f39", x"7f39", x"7f39", x"7f38", x"7f38", x"7f38", 
    x"7f37", x"7f37", x"7f37", x"7f36", x"7f36", x"7f36", x"7f35", x"7f35", 
    x"7f35", x"7f34", x"7f34", x"7f34", x"7f33", x"7f33", x"7f32", x"7f32", 
    x"7f32", x"7f31", x"7f31", x"7f31", x"7f30", x"7f30", x"7f30", x"7f2f", 
    x"7f2f", x"7f2f", x"7f2e", x"7f2e", x"7f2e", x"7f2d", x"7f2d", x"7f2c", 
    x"7f2c", x"7f2c", x"7f2b", x"7f2b", x"7f2b", x"7f2a", x"7f2a", x"7f2a", 
    x"7f29", x"7f29", x"7f29", x"7f28", x"7f28", x"7f27", x"7f27", x"7f27", 
    x"7f26", x"7f26", x"7f26", x"7f25", x"7f25", x"7f25", x"7f24", x"7f24", 
    x"7f23", x"7f23", x"7f23", x"7f22", x"7f22", x"7f22", x"7f21", x"7f21", 
    x"7f21", x"7f20", x"7f20", x"7f1f", x"7f1f", x"7f1f", x"7f1e", x"7f1e", 
    x"7f1e", x"7f1d", x"7f1d", x"7f1d", x"7f1c", x"7f1c", x"7f1b", x"7f1b", 
    x"7f1b", x"7f1a", x"7f1a", x"7f1a", x"7f19", x"7f19", x"7f18", x"7f18", 
    x"7f18", x"7f17", x"7f17", x"7f17", x"7f16", x"7f16", x"7f15", x"7f15", 
    x"7f15", x"7f14", x"7f14", x"7f14", x"7f13", x"7f13", x"7f12", x"7f12", 
    x"7f12", x"7f11", x"7f11", x"7f11", x"7f10", x"7f10", x"7f0f", x"7f0f", 
    x"7f0f", x"7f0e", x"7f0e", x"7f0e", x"7f0d", x"7f0d", x"7f0c", x"7f0c", 
    x"7f0c", x"7f0b", x"7f0b", x"7f0a", x"7f0a", x"7f0a", x"7f09", x"7f09", 
    x"7f09", x"7f08", x"7f08", x"7f07", x"7f07", x"7f07", x"7f06", x"7f06", 
    x"7f05", x"7f05", x"7f05", x"7f04", x"7f04", x"7f04", x"7f03", x"7f03", 
    x"7f02", x"7f02", x"7f02", x"7f01", x"7f01", x"7f00", x"7f00", x"7f00", 
    x"7eff", x"7eff", x"7efe", x"7efe", x"7efe", x"7efd", x"7efd", x"7efd", 
    x"7efc", x"7efc", x"7efb", x"7efb", x"7efb", x"7efa", x"7efa", x"7ef9", 
    x"7ef9", x"7ef9", x"7ef8", x"7ef8", x"7ef7", x"7ef7", x"7ef7", x"7ef6", 
    x"7ef6", x"7ef5", x"7ef5", x"7ef5", x"7ef4", x"7ef4", x"7ef3", x"7ef3", 
    x"7ef3", x"7ef2", x"7ef2", x"7ef1", x"7ef1", x"7ef1", x"7ef0", x"7ef0", 
    x"7eef", x"7eef", x"7eef", x"7eee", x"7eee", x"7eed", x"7eed", x"7eed", 
    x"7eec", x"7eec", x"7eeb", x"7eeb", x"7eea", x"7eea", x"7eea", x"7ee9", 
    x"7ee9", x"7ee8", x"7ee8", x"7ee8", x"7ee7", x"7ee7", x"7ee6", x"7ee6", 
    x"7ee6", x"7ee5", x"7ee5", x"7ee4", x"7ee4", x"7ee4", x"7ee3", x"7ee3", 
    x"7ee2", x"7ee2", x"7ee1", x"7ee1", x"7ee1", x"7ee0", x"7ee0", x"7edf", 
    x"7edf", x"7edf", x"7ede", x"7ede", x"7edd", x"7edd", x"7edc", x"7edc", 
    x"7edc", x"7edb", x"7edb", x"7eda", x"7eda", x"7eda", x"7ed9", x"7ed9", 
    x"7ed8", x"7ed8", x"7ed7", x"7ed7", x"7ed7", x"7ed6", x"7ed6", x"7ed5", 
    x"7ed5", x"7ed4", x"7ed4", x"7ed4", x"7ed3", x"7ed3", x"7ed2", x"7ed2", 
    x"7ed2", x"7ed1", x"7ed1", x"7ed0", x"7ed0", x"7ecf", x"7ecf", x"7ecf", 
    x"7ece", x"7ece", x"7ecd", x"7ecd", x"7ecc", x"7ecc", x"7ecc", x"7ecb", 
    x"7ecb", x"7eca", x"7eca", x"7ec9", x"7ec9", x"7ec9", x"7ec8", x"7ec8", 
    x"7ec7", x"7ec7", x"7ec6", x"7ec6", x"7ec5", x"7ec5", x"7ec5", x"7ec4", 
    x"7ec4", x"7ec3", x"7ec3", x"7ec2", x"7ec2", x"7ec2", x"7ec1", x"7ec1", 
    x"7ec0", x"7ec0", x"7ebf", x"7ebf", x"7ebf", x"7ebe", x"7ebe", x"7ebd", 
    x"7ebd", x"7ebc", x"7ebc", x"7ebb", x"7ebb", x"7ebb", x"7eba", x"7eba", 
    x"7eb9", x"7eb9", x"7eb8", x"7eb8", x"7eb7", x"7eb7", x"7eb7", x"7eb6", 
    x"7eb6", x"7eb5", x"7eb5", x"7eb4", x"7eb4", x"7eb3", x"7eb3", x"7eb3", 
    x"7eb2", x"7eb2", x"7eb1", x"7eb1", x"7eb0", x"7eb0", x"7eaf", x"7eaf", 
    x"7eaf", x"7eae", x"7eae", x"7ead", x"7ead", x"7eac", x"7eac", x"7eab", 
    x"7eab", x"7eaa", x"7eaa", x"7eaa", x"7ea9", x"7ea9", x"7ea8", x"7ea8", 
    x"7ea7", x"7ea7", x"7ea6", x"7ea6", x"7ea6", x"7ea5", x"7ea5", x"7ea4", 
    x"7ea4", x"7ea3", x"7ea3", x"7ea2", x"7ea2", x"7ea1", x"7ea1", x"7ea0", 
    x"7ea0", x"7ea0", x"7e9f", x"7e9f", x"7e9e", x"7e9e", x"7e9d", x"7e9d", 
    x"7e9c", x"7e9c", x"7e9b", x"7e9b", x"7e9b", x"7e9a", x"7e9a", x"7e99", 
    x"7e99", x"7e98", x"7e98", x"7e97", x"7e97", x"7e96", x"7e96", x"7e95", 
    x"7e95", x"7e94", x"7e94", x"7e94", x"7e93", x"7e93", x"7e92", x"7e92", 
    x"7e91", x"7e91", x"7e90", x"7e90", x"7e8f", x"7e8f", x"7e8e", x"7e8e", 
    x"7e8d", x"7e8d", x"7e8d", x"7e8c", x"7e8c", x"7e8b", x"7e8b", x"7e8a", 
    x"7e8a", x"7e89", x"7e89", x"7e88", x"7e88", x"7e87", x"7e87", x"7e86", 
    x"7e86", x"7e85", x"7e85", x"7e84", x"7e84", x"7e83", x"7e83", x"7e83", 
    x"7e82", x"7e82", x"7e81", x"7e81", x"7e80", x"7e80", x"7e7f", x"7e7f", 
    x"7e7e", x"7e7e", x"7e7d", x"7e7d", x"7e7c", x"7e7c", x"7e7b", x"7e7b", 
    x"7e7a", x"7e7a", x"7e79", x"7e79", x"7e78", x"7e78", x"7e77", x"7e77", 
    x"7e77", x"7e76", x"7e76", x"7e75", x"7e75", x"7e74", x"7e74", x"7e73", 
    x"7e73", x"7e72", x"7e72", x"7e71", x"7e71", x"7e70", x"7e70", x"7e6f", 
    x"7e6f", x"7e6e", x"7e6e", x"7e6d", x"7e6d", x"7e6c", x"7e6c", x"7e6b", 
    x"7e6b", x"7e6a", x"7e6a", x"7e69", x"7e69", x"7e68", x"7e68", x"7e67", 
    x"7e67", x"7e66", x"7e66", x"7e65", x"7e65", x"7e64", x"7e64", x"7e63", 
    x"7e63", x"7e62", x"7e62", x"7e61", x"7e61", x"7e60", x"7e60", x"7e5f", 
    x"7e5f", x"7e5e", x"7e5e", x"7e5d", x"7e5d", x"7e5c", x"7e5c", x"7e5b", 
    x"7e5b", x"7e5a", x"7e5a", x"7e59", x"7e59", x"7e58", x"7e58", x"7e57", 
    x"7e57", x"7e56", x"7e56", x"7e55", x"7e55", x"7e54", x"7e54", x"7e53", 
    x"7e53", x"7e52", x"7e52", x"7e51", x"7e51", x"7e50", x"7e50", x"7e4f", 
    x"7e4f", x"7e4e", x"7e4e", x"7e4d", x"7e4d", x"7e4c", x"7e4c", x"7e4b", 
    x"7e4b", x"7e4a", x"7e4a", x"7e49", x"7e49", x"7e48", x"7e48", x"7e47", 
    x"7e47", x"7e46", x"7e46", x"7e45", x"7e45", x"7e44", x"7e44", x"7e43", 
    x"7e42", x"7e42", x"7e41", x"7e41", x"7e40", x"7e40", x"7e3f", x"7e3f", 
    x"7e3e", x"7e3e", x"7e3d", x"7e3d", x"7e3c", x"7e3c", x"7e3b", x"7e3b", 
    x"7e3a", x"7e3a", x"7e39", x"7e39", x"7e38", x"7e38", x"7e37", x"7e37", 
    x"7e36", x"7e36", x"7e35", x"7e34", x"7e34", x"7e33", x"7e33", x"7e32", 
    x"7e32", x"7e31", x"7e31", x"7e30", x"7e30", x"7e2f", x"7e2f", x"7e2e", 
    x"7e2e", x"7e2d", x"7e2d", x"7e2c", x"7e2c", x"7e2b", x"7e2a", x"7e2a", 
    x"7e29", x"7e29", x"7e28", x"7e28", x"7e27", x"7e27", x"7e26", x"7e26", 
    x"7e25", x"7e25", x"7e24", x"7e24", x"7e23", x"7e22", x"7e22", x"7e21", 
    x"7e21", x"7e20", x"7e20", x"7e1f", x"7e1f", x"7e1e", x"7e1e", x"7e1d", 
    x"7e1d", x"7e1c", x"7e1c", x"7e1b", x"7e1a", x"7e1a", x"7e19", x"7e19", 
    x"7e18", x"7e18", x"7e17", x"7e17", x"7e16", x"7e16", x"7e15", x"7e15", 
    x"7e14", x"7e13", x"7e13", x"7e12", x"7e12", x"7e11", x"7e11", x"7e10", 
    x"7e10", x"7e0f", x"7e0f", x"7e0e", x"7e0d", x"7e0d", x"7e0c", x"7e0c", 
    x"7e0b", x"7e0b", x"7e0a", x"7e0a", x"7e09", x"7e09", x"7e08", x"7e07", 
    x"7e07", x"7e06", x"7e06", x"7e05", x"7e05", x"7e04", x"7e04", x"7e03", 
    x"7e02", x"7e02", x"7e01", x"7e01", x"7e00", x"7e00", x"7dff", x"7dff", 
    x"7dfe", x"7dfd", x"7dfd", x"7dfc", x"7dfc", x"7dfb", x"7dfb", x"7dfa", 
    x"7dfa", x"7df9", x"7df8", x"7df8", x"7df7", x"7df7", x"7df6", x"7df6", 
    x"7df5", x"7df5", x"7df4", x"7df3", x"7df3", x"7df2", x"7df2", x"7df1", 
    x"7df1", x"7df0", x"7df0", x"7def", x"7dee", x"7dee", x"7ded", x"7ded", 
    x"7dec", x"7dec", x"7deb", x"7dea", x"7dea", x"7de9", x"7de9", x"7de8", 
    x"7de8", x"7de7", x"7de7", x"7de6", x"7de5", x"7de5", x"7de4", x"7de4", 
    x"7de3", x"7de3", x"7de2", x"7de1", x"7de1", x"7de0", x"7de0", x"7ddf", 
    x"7ddf", x"7dde", x"7ddd", x"7ddd", x"7ddc", x"7ddc", x"7ddb", x"7ddb", 
    x"7dda", x"7dd9", x"7dd9", x"7dd8", x"7dd8", x"7dd7", x"7dd7", x"7dd6", 
    x"7dd5", x"7dd5", x"7dd4", x"7dd4", x"7dd3", x"7dd3", x"7dd2", x"7dd1", 
    x"7dd1", x"7dd0", x"7dd0", x"7dcf", x"7dce", x"7dce", x"7dcd", x"7dcd", 
    x"7dcc", x"7dcc", x"7dcb", x"7dca", x"7dca", x"7dc9", x"7dc9", x"7dc8", 
    x"7dc8", x"7dc7", x"7dc6", x"7dc6", x"7dc5", x"7dc5", x"7dc4", x"7dc3", 
    x"7dc3", x"7dc2", x"7dc2", x"7dc1", x"7dc1", x"7dc0", x"7dbf", x"7dbf", 
    x"7dbe", x"7dbe", x"7dbd", x"7dbc", x"7dbc", x"7dbb", x"7dbb", x"7dba", 
    x"7db9", x"7db9", x"7db8", x"7db8", x"7db7", x"7db7", x"7db6", x"7db5", 
    x"7db5", x"7db4", x"7db4", x"7db3", x"7db2", x"7db2", x"7db1", x"7db1", 
    x"7db0", x"7daf", x"7daf", x"7dae", x"7dae", x"7dad", x"7dac", x"7dac", 
    x"7dab", x"7dab", x"7daa", x"7da9", x"7da9", x"7da8", x"7da8", x"7da7", 
    x"7da6", x"7da6", x"7da5", x"7da5", x"7da4", x"7da3", x"7da3", x"7da2", 
    x"7da2", x"7da1", x"7da0", x"7da0", x"7d9f", x"7d9f", x"7d9e", x"7d9d", 
    x"7d9d", x"7d9c", x"7d9c", x"7d9b", x"7d9a", x"7d9a", x"7d99", x"7d99", 
    x"7d98", x"7d97", x"7d97", x"7d96", x"7d96", x"7d95", x"7d94", x"7d94", 
    x"7d93", x"7d93", x"7d92", x"7d91", x"7d91", x"7d90", x"7d90", x"7d8f", 
    x"7d8e", x"7d8e", x"7d8d", x"7d8c", x"7d8c", x"7d8b", x"7d8b", x"7d8a", 
    x"7d89", x"7d89", x"7d88", x"7d88", x"7d87", x"7d86", x"7d86", x"7d85", 
    x"7d84", x"7d84", x"7d83", x"7d83", x"7d82", x"7d81", x"7d81", x"7d80", 
    x"7d80", x"7d7f", x"7d7e", x"7d7e", x"7d7d", x"7d7c", x"7d7c", x"7d7b", 
    x"7d7b", x"7d7a", x"7d79", x"7d79", x"7d78", x"7d77", x"7d77", x"7d76", 
    x"7d76", x"7d75", x"7d74", x"7d74", x"7d73", x"7d73", x"7d72", x"7d71", 
    x"7d71", x"7d70", x"7d6f", x"7d6f", x"7d6e", x"7d6e", x"7d6d", x"7d6c", 
    x"7d6c", x"7d6b", x"7d6a", x"7d6a", x"7d69", x"7d68", x"7d68", x"7d67", 
    x"7d67", x"7d66", x"7d65", x"7d65", x"7d64", x"7d63", x"7d63", x"7d62", 
    x"7d62", x"7d61", x"7d60", x"7d60", x"7d5f", x"7d5e", x"7d5e", x"7d5d", 
    x"7d5c", x"7d5c", x"7d5b", x"7d5b", x"7d5a", x"7d59", x"7d59", x"7d58", 
    x"7d57", x"7d57", x"7d56", x"7d56", x"7d55", x"7d54", x"7d54", x"7d53", 
    x"7d52", x"7d52", x"7d51", x"7d50", x"7d50", x"7d4f", x"7d4e", x"7d4e", 
    x"7d4d", x"7d4d", x"7d4c", x"7d4b", x"7d4b", x"7d4a", x"7d49", x"7d49", 
    x"7d48", x"7d47", x"7d47", x"7d46", x"7d45", x"7d45", x"7d44", x"7d44", 
    x"7d43", x"7d42", x"7d42", x"7d41", x"7d40", x"7d40", x"7d3f", x"7d3e", 
    x"7d3e", x"7d3d", x"7d3c", x"7d3c", x"7d3b", x"7d3a", x"7d3a", x"7d39", 
    x"7d39", x"7d38", x"7d37", x"7d37", x"7d36", x"7d35", x"7d35", x"7d34", 
    x"7d33", x"7d33", x"7d32", x"7d31", x"7d31", x"7d30", x"7d2f", x"7d2f", 
    x"7d2e", x"7d2d", x"7d2d", x"7d2c", x"7d2b", x"7d2b", x"7d2a", x"7d29", 
    x"7d29", x"7d28", x"7d28", x"7d27", x"7d26", x"7d26", x"7d25", x"7d24", 
    x"7d24", x"7d23", x"7d22", x"7d22", x"7d21", x"7d20", x"7d20", x"7d1f", 
    x"7d1e", x"7d1e", x"7d1d", x"7d1c", x"7d1c", x"7d1b", x"7d1a", x"7d1a", 
    x"7d19", x"7d18", x"7d18", x"7d17", x"7d16", x"7d16", x"7d15", x"7d14", 
    x"7d14", x"7d13", x"7d12", x"7d12", x"7d11", x"7d10", x"7d10", x"7d0f", 
    x"7d0e", x"7d0e", x"7d0d", x"7d0c", x"7d0c", x"7d0b", x"7d0a", x"7d0a", 
    x"7d09", x"7d08", x"7d08", x"7d07", x"7d06", x"7d06", x"7d05", x"7d04", 
    x"7d04", x"7d03", x"7d02", x"7d02", x"7d01", x"7d00", x"7cff", x"7cff", 
    x"7cfe", x"7cfd", x"7cfd", x"7cfc", x"7cfb", x"7cfb", x"7cfa", x"7cf9", 
    x"7cf9", x"7cf8", x"7cf7", x"7cf7", x"7cf6", x"7cf5", x"7cf5", x"7cf4", 
    x"7cf3", x"7cf3", x"7cf2", x"7cf1", x"7cf1", x"7cf0", x"7cef", x"7cee", 
    x"7cee", x"7ced", x"7cec", x"7cec", x"7ceb", x"7cea", x"7cea", x"7ce9", 
    x"7ce8", x"7ce8", x"7ce7", x"7ce6", x"7ce6", x"7ce5", x"7ce4", x"7ce4", 
    x"7ce3", x"7ce2", x"7ce1", x"7ce1", x"7ce0", x"7cdf", x"7cdf", x"7cde", 
    x"7cdd", x"7cdd", x"7cdc", x"7cdb", x"7cdb", x"7cda", x"7cd9", x"7cd8", 
    x"7cd8", x"7cd7", x"7cd6", x"7cd6", x"7cd5", x"7cd4", x"7cd4", x"7cd3", 
    x"7cd2", x"7cd2", x"7cd1", x"7cd0", x"7ccf", x"7ccf", x"7cce", x"7ccd", 
    x"7ccd", x"7ccc", x"7ccb", x"7ccb", x"7cca", x"7cc9", x"7cc8", x"7cc8", 
    x"7cc7", x"7cc6", x"7cc6", x"7cc5", x"7cc4", x"7cc4", x"7cc3", x"7cc2", 
    x"7cc1", x"7cc1", x"7cc0", x"7cbf", x"7cbf", x"7cbe", x"7cbd", x"7cbd", 
    x"7cbc", x"7cbb", x"7cba", x"7cba", x"7cb9", x"7cb8", x"7cb8", x"7cb7", 
    x"7cb6", x"7cb5", x"7cb5", x"7cb4", x"7cb3", x"7cb3", x"7cb2", x"7cb1", 
    x"7cb1", x"7cb0", x"7caf", x"7cae", x"7cae", x"7cad", x"7cac", x"7cac", 
    x"7cab", x"7caa", x"7ca9", x"7ca9", x"7ca8", x"7ca7", x"7ca7", x"7ca6", 
    x"7ca5", x"7ca4", x"7ca4", x"7ca3", x"7ca2", x"7ca2", x"7ca1", x"7ca0", 
    x"7c9f", x"7c9f", x"7c9e", x"7c9d", x"7c9d", x"7c9c", x"7c9b", x"7c9a", 
    x"7c9a", x"7c99", x"7c98", x"7c98", x"7c97", x"7c96", x"7c95", x"7c95", 
    x"7c94", x"7c93", x"7c92", x"7c92", x"7c91", x"7c90", x"7c90", x"7c8f", 
    x"7c8e", x"7c8d", x"7c8d", x"7c8c", x"7c8b", x"7c8a", x"7c8a", x"7c89", 
    x"7c88", x"7c88", x"7c87", x"7c86", x"7c85", x"7c85", x"7c84", x"7c83", 
    x"7c83", x"7c82", x"7c81", x"7c80", x"7c80", x"7c7f", x"7c7e", x"7c7d", 
    x"7c7d", x"7c7c", x"7c7b", x"7c7a", x"7c7a", x"7c79", x"7c78", x"7c78", 
    x"7c77", x"7c76", x"7c75", x"7c75", x"7c74", x"7c73", x"7c72", x"7c72", 
    x"7c71", x"7c70", x"7c6f", x"7c6f", x"7c6e", x"7c6d", x"7c6d", x"7c6c", 
    x"7c6b", x"7c6a", x"7c6a", x"7c69", x"7c68", x"7c67", x"7c67", x"7c66", 
    x"7c65", x"7c64", x"7c64", x"7c63", x"7c62", x"7c61", x"7c61", x"7c60", 
    x"7c5f", x"7c5e", x"7c5e", x"7c5d", x"7c5c", x"7c5c", x"7c5b", x"7c5a", 
    x"7c59", x"7c59", x"7c58", x"7c57", x"7c56", x"7c56", x"7c55", x"7c54", 
    x"7c53", x"7c53", x"7c52", x"7c51", x"7c50", x"7c50", x"7c4f", x"7c4e", 
    x"7c4d", x"7c4d", x"7c4c", x"7c4b", x"7c4a", x"7c4a", x"7c49", x"7c48", 
    x"7c47", x"7c47", x"7c46", x"7c45", x"7c44", x"7c44", x"7c43", x"7c42", 
    x"7c41", x"7c41", x"7c40", x"7c3f", x"7c3e", x"7c3e", x"7c3d", x"7c3c", 
    x"7c3b", x"7c3a", x"7c3a", x"7c39", x"7c38", x"7c37", x"7c37", x"7c36", 
    x"7c35", x"7c34", x"7c34", x"7c33", x"7c32", x"7c31", x"7c31", x"7c30", 
    x"7c2f", x"7c2e", x"7c2e", x"7c2d", x"7c2c", x"7c2b", x"7c2b", x"7c2a", 
    x"7c29", x"7c28", x"7c27", x"7c27", x"7c26", x"7c25", x"7c24", x"7c24", 
    x"7c23", x"7c22", x"7c21", x"7c21", x"7c20", x"7c1f", x"7c1e", x"7c1e", 
    x"7c1d", x"7c1c", x"7c1b", x"7c1a", x"7c1a", x"7c19", x"7c18", x"7c17", 
    x"7c17", x"7c16", x"7c15", x"7c14", x"7c14", x"7c13", x"7c12", x"7c11", 
    x"7c10", x"7c10", x"7c0f", x"7c0e", x"7c0d", x"7c0d", x"7c0c", x"7c0b", 
    x"7c0a", x"7c09", x"7c09", x"7c08", x"7c07", x"7c06", x"7c06", x"7c05", 
    x"7c04", x"7c03", x"7c02", x"7c02", x"7c01", x"7c00", x"7bff", x"7bff", 
    x"7bfe", x"7bfd", x"7bfc", x"7bfb", x"7bfb", x"7bfa", x"7bf9", x"7bf8", 
    x"7bf8", x"7bf7", x"7bf6", x"7bf5", x"7bf4", x"7bf4", x"7bf3", x"7bf2", 
    x"7bf1", x"7bf1", x"7bf0", x"7bef", x"7bee", x"7bed", x"7bed", x"7bec", 
    x"7beb", x"7bea", x"7be9", x"7be9", x"7be8", x"7be7", x"7be6", x"7be6", 
    x"7be5", x"7be4", x"7be3", x"7be2", x"7be2", x"7be1", x"7be0", x"7bdf", 
    x"7bde", x"7bde", x"7bdd", x"7bdc", x"7bdb", x"7bda", x"7bda", x"7bd9", 
    x"7bd8", x"7bd7", x"7bd6", x"7bd6", x"7bd5", x"7bd4", x"7bd3", x"7bd2", 
    x"7bd2", x"7bd1", x"7bd0", x"7bcf", x"7bcf", x"7bce", x"7bcd", x"7bcc", 
    x"7bcb", x"7bcb", x"7bca", x"7bc9", x"7bc8", x"7bc7", x"7bc7", x"7bc6", 
    x"7bc5", x"7bc4", x"7bc3", x"7bc3", x"7bc2", x"7bc1", x"7bc0", x"7bbf", 
    x"7bbf", x"7bbe", x"7bbd", x"7bbc", x"7bbb", x"7bba", x"7bba", x"7bb9", 
    x"7bb8", x"7bb7", x"7bb6", x"7bb6", x"7bb5", x"7bb4", x"7bb3", x"7bb2", 
    x"7bb2", x"7bb1", x"7bb0", x"7baf", x"7bae", x"7bae", x"7bad", x"7bac", 
    x"7bab", x"7baa", x"7baa", x"7ba9", x"7ba8", x"7ba7", x"7ba6", x"7ba5", 
    x"7ba5", x"7ba4", x"7ba3", x"7ba2", x"7ba1", x"7ba1", x"7ba0", x"7b9f", 
    x"7b9e", x"7b9d", x"7b9d", x"7b9c", x"7b9b", x"7b9a", x"7b99", x"7b98", 
    x"7b98", x"7b97", x"7b96", x"7b95", x"7b94", x"7b94", x"7b93", x"7b92", 
    x"7b91", x"7b90", x"7b8f", x"7b8f", x"7b8e", x"7b8d", x"7b8c", x"7b8b", 
    x"7b8b", x"7b8a", x"7b89", x"7b88", x"7b87", x"7b86", x"7b86", x"7b85", 
    x"7b84", x"7b83", x"7b82", x"7b81", x"7b81", x"7b80", x"7b7f", x"7b7e", 
    x"7b7d", x"7b7d", x"7b7c", x"7b7b", x"7b7a", x"7b79", x"7b78", x"7b78", 
    x"7b77", x"7b76", x"7b75", x"7b74", x"7b73", x"7b73", x"7b72", x"7b71", 
    x"7b70", x"7b6f", x"7b6e", x"7b6e", x"7b6d", x"7b6c", x"7b6b", x"7b6a", 
    x"7b69", x"7b69", x"7b68", x"7b67", x"7b66", x"7b65", x"7b64", x"7b64", 
    x"7b63", x"7b62", x"7b61", x"7b60", x"7b5f", x"7b5f", x"7b5e", x"7b5d", 
    x"7b5c", x"7b5b", x"7b5a", x"7b5a", x"7b59", x"7b58", x"7b57", x"7b56", 
    x"7b55", x"7b54", x"7b54", x"7b53", x"7b52", x"7b51", x"7b50", x"7b4f", 
    x"7b4f", x"7b4e", x"7b4d", x"7b4c", x"7b4b", x"7b4a", x"7b4a", x"7b49", 
    x"7b48", x"7b47", x"7b46", x"7b45", x"7b44", x"7b44", x"7b43", x"7b42", 
    x"7b41", x"7b40", x"7b3f", x"7b3f", x"7b3e", x"7b3d", x"7b3c", x"7b3b", 
    x"7b3a", x"7b39", x"7b39", x"7b38", x"7b37", x"7b36", x"7b35", x"7b34", 
    x"7b33", x"7b33", x"7b32", x"7b31", x"7b30", x"7b2f", x"7b2e", x"7b2e", 
    x"7b2d", x"7b2c", x"7b2b", x"7b2a", x"7b29", x"7b28", x"7b28", x"7b27", 
    x"7b26", x"7b25", x"7b24", x"7b23", x"7b22", x"7b22", x"7b21", x"7b20", 
    x"7b1f", x"7b1e", x"7b1d", x"7b1c", x"7b1c", x"7b1b", x"7b1a", x"7b19", 
    x"7b18", x"7b17", x"7b16", x"7b16", x"7b15", x"7b14", x"7b13", x"7b12", 
    x"7b11", x"7b10", x"7b0f", x"7b0f", x"7b0e", x"7b0d", x"7b0c", x"7b0b", 
    x"7b0a", x"7b09", x"7b09", x"7b08", x"7b07", x"7b06", x"7b05", x"7b04", 
    x"7b03", x"7b02", x"7b02", x"7b01", x"7b00", x"7aff", x"7afe", x"7afd", 
    x"7afc", x"7afc", x"7afb", x"7afa", x"7af9", x"7af8", x"7af7", x"7af6", 
    x"7af5", x"7af5", x"7af4", x"7af3", x"7af2", x"7af1", x"7af0", x"7aef", 
    x"7aee", x"7aee", x"7aed", x"7aec", x"7aeb", x"7aea", x"7ae9", x"7ae8", 
    x"7ae7", x"7ae7", x"7ae6", x"7ae5", x"7ae4", x"7ae3", x"7ae2", x"7ae1", 
    x"7ae0", x"7ae0", x"7adf", x"7ade", x"7add", x"7adc", x"7adb", x"7ada", 
    x"7ad9", x"7ad8", x"7ad8", x"7ad7", x"7ad6", x"7ad5", x"7ad4", x"7ad3", 
    x"7ad2", x"7ad1", x"7ad1", x"7ad0", x"7acf", x"7ace", x"7acd", x"7acc", 
    x"7acb", x"7aca", x"7ac9", x"7ac9", x"7ac8", x"7ac7", x"7ac6", x"7ac5", 
    x"7ac4", x"7ac3", x"7ac2", x"7ac1", x"7ac1", x"7ac0", x"7abf", x"7abe", 
    x"7abd", x"7abc", x"7abb", x"7aba", x"7ab9", x"7ab9", x"7ab8", x"7ab7", 
    x"7ab6", x"7ab5", x"7ab4", x"7ab3", x"7ab2", x"7ab1", x"7ab0", x"7ab0", 
    x"7aaf", x"7aae", x"7aad", x"7aac", x"7aab", x"7aaa", x"7aa9", x"7aa8", 
    x"7aa8", x"7aa7", x"7aa6", x"7aa5", x"7aa4", x"7aa3", x"7aa2", x"7aa1", 
    x"7aa0", x"7a9f", x"7a9f", x"7a9e", x"7a9d", x"7a9c", x"7a9b", x"7a9a", 
    x"7a99", x"7a98", x"7a97", x"7a96", x"7a95", x"7a95", x"7a94", x"7a93", 
    x"7a92", x"7a91", x"7a90", x"7a8f", x"7a8e", x"7a8d", x"7a8c", x"7a8c", 
    x"7a8b", x"7a8a", x"7a89", x"7a88", x"7a87", x"7a86", x"7a85", x"7a84", 
    x"7a83", x"7a82", x"7a82", x"7a81", x"7a80", x"7a7f", x"7a7e", x"7a7d", 
    x"7a7c", x"7a7b", x"7a7a", x"7a79", x"7a78", x"7a78", x"7a77", x"7a76", 
    x"7a75", x"7a74", x"7a73", x"7a72", x"7a71", x"7a70", x"7a6f", x"7a6e", 
    x"7a6d", x"7a6d", x"7a6c", x"7a6b", x"7a6a", x"7a69", x"7a68", x"7a67", 
    x"7a66", x"7a65", x"7a64", x"7a63", x"7a62", x"7a61", x"7a61", x"7a60", 
    x"7a5f", x"7a5e", x"7a5d", x"7a5c", x"7a5b", x"7a5a", x"7a59", x"7a58", 
    x"7a57", x"7a56", x"7a56", x"7a55", x"7a54", x"7a53", x"7a52", x"7a51", 
    x"7a50", x"7a4f", x"7a4e", x"7a4d", x"7a4c", x"7a4b", x"7a4a", x"7a49", 
    x"7a49", x"7a48", x"7a47", x"7a46", x"7a45", x"7a44", x"7a43", x"7a42", 
    x"7a41", x"7a40", x"7a3f", x"7a3e", x"7a3d", x"7a3c", x"7a3c", x"7a3b", 
    x"7a3a", x"7a39", x"7a38", x"7a37", x"7a36", x"7a35", x"7a34", x"7a33", 
    x"7a32", x"7a31", x"7a30", x"7a2f", x"7a2e", x"7a2e", x"7a2d", x"7a2c", 
    x"7a2b", x"7a2a", x"7a29", x"7a28", x"7a27", x"7a26", x"7a25", x"7a24", 
    x"7a23", x"7a22", x"7a21", x"7a20", x"7a1f", x"7a1e", x"7a1e", x"7a1d", 
    x"7a1c", x"7a1b", x"7a1a", x"7a19", x"7a18", x"7a17", x"7a16", x"7a15", 
    x"7a14", x"7a13", x"7a12", x"7a11", x"7a10", x"7a0f", x"7a0e", x"7a0e", 
    x"7a0d", x"7a0c", x"7a0b", x"7a0a", x"7a09", x"7a08", x"7a07", x"7a06", 
    x"7a05", x"7a04", x"7a03", x"7a02", x"7a01", x"7a00", x"79ff", x"79fe", 
    x"79fd", x"79fc", x"79fb", x"79fb", x"79fa", x"79f9", x"79f8", x"79f7", 
    x"79f6", x"79f5", x"79f4", x"79f3", x"79f2", x"79f1", x"79f0", x"79ef", 
    x"79ee", x"79ed", x"79ec", x"79eb", x"79ea", x"79e9", x"79e8", x"79e7", 
    x"79e6", x"79e6", x"79e5", x"79e4", x"79e3", x"79e2", x"79e1", x"79e0", 
    x"79df", x"79de", x"79dd", x"79dc", x"79db", x"79da", x"79d9", x"79d8", 
    x"79d7", x"79d6", x"79d5", x"79d4", x"79d3", x"79d2", x"79d1", x"79d0", 
    x"79cf", x"79ce", x"79cd", x"79cd", x"79cc", x"79cb", x"79ca", x"79c9", 
    x"79c8", x"79c7", x"79c6", x"79c5", x"79c4", x"79c3", x"79c2", x"79c1", 
    x"79c0", x"79bf", x"79be", x"79bd", x"79bc", x"79bb", x"79ba", x"79b9", 
    x"79b8", x"79b7", x"79b6", x"79b5", x"79b4", x"79b3", x"79b2", x"79b1", 
    x"79b0", x"79af", x"79ae", x"79ad", x"79ac", x"79ac", x"79ab", x"79aa", 
    x"79a9", x"79a8", x"79a7", x"79a6", x"79a5", x"79a4", x"79a3", x"79a2", 
    x"79a1", x"79a0", x"799f", x"799e", x"799d", x"799c", x"799b", x"799a", 
    x"7999", x"7998", x"7997", x"7996", x"7995", x"7994", x"7993", x"7992", 
    x"7991", x"7990", x"798f", x"798e", x"798d", x"798c", x"798b", x"798a", 
    x"7989", x"7988", x"7987", x"7986", x"7985", x"7984", x"7983", x"7982", 
    x"7981", x"7980", x"797f", x"797e", x"797d", x"797c", x"797b", x"797a", 
    x"7979", x"7978", x"7977", x"7976", x"7975", x"7974", x"7973", x"7972", 
    x"7971", x"7970", x"796f", x"796e", x"796d", x"796c", x"796b", x"796b", 
    x"796a", x"7969", x"7968", x"7967", x"7966", x"7965", x"7964", x"7963", 
    x"7962", x"7961", x"7960", x"795f", x"795e", x"795d", x"795c", x"795b", 
    x"795a", x"7959", x"7958", x"7957", x"7956", x"7955", x"7954", x"7953", 
    x"7952", x"7951", x"7950", x"794f", x"794e", x"794d", x"794c", x"794b", 
    x"794a", x"7949", x"7948", x"7947", x"7946", x"7945", x"7944", x"7943", 
    x"7941", x"7940", x"793f", x"793e", x"793d", x"793c", x"793b", x"793a", 
    x"7939", x"7938", x"7937", x"7936", x"7935", x"7934", x"7933", x"7932", 
    x"7931", x"7930", x"792f", x"792e", x"792d", x"792c", x"792b", x"792a", 
    x"7929", x"7928", x"7927", x"7926", x"7925", x"7924", x"7923", x"7922", 
    x"7921", x"7920", x"791f", x"791e", x"791d", x"791c", x"791b", x"791a", 
    x"7919", x"7918", x"7917", x"7916", x"7915", x"7914", x"7913", x"7912", 
    x"7911", x"7910", x"790f", x"790e", x"790d", x"790c", x"790b", x"790a", 
    x"7909", x"7908", x"7907", x"7906", x"7905", x"7904", x"7903", x"7902", 
    x"7901", x"7900", x"78fe", x"78fd", x"78fc", x"78fb", x"78fa", x"78f9", 
    x"78f8", x"78f7", x"78f6", x"78f5", x"78f4", x"78f3", x"78f2", x"78f1", 
    x"78f0", x"78ef", x"78ee", x"78ed", x"78ec", x"78eb", x"78ea", x"78e9", 
    x"78e8", x"78e7", x"78e6", x"78e5", x"78e4", x"78e3", x"78e2", x"78e1", 
    x"78e0", x"78df", x"78de", x"78dd", x"78db", x"78da", x"78d9", x"78d8", 
    x"78d7", x"78d6", x"78d5", x"78d4", x"78d3", x"78d2", x"78d1", x"78d0", 
    x"78cf", x"78ce", x"78cd", x"78cc", x"78cb", x"78ca", x"78c9", x"78c8", 
    x"78c7", x"78c6", x"78c5", x"78c4", x"78c3", x"78c2", x"78c0", x"78bf", 
    x"78be", x"78bd", x"78bc", x"78bb", x"78ba", x"78b9", x"78b8", x"78b7", 
    x"78b6", x"78b5", x"78b4", x"78b3", x"78b2", x"78b1", x"78b0", x"78af", 
    x"78ae", x"78ad", x"78ac", x"78ab", x"78a9", x"78a8", x"78a7", x"78a6", 
    x"78a5", x"78a4", x"78a3", x"78a2", x"78a1", x"78a0", x"789f", x"789e", 
    x"789d", x"789c", x"789b", x"789a", x"7899", x"7898", x"7897", x"7896", 
    x"7894", x"7893", x"7892", x"7891", x"7890", x"788f", x"788e", x"788d", 
    x"788c", x"788b", x"788a", x"7889", x"7888", x"7887", x"7886", x"7885", 
    x"7884", x"7883", x"7881", x"7880", x"787f", x"787e", x"787d", x"787c", 
    x"787b", x"787a", x"7879", x"7878", x"7877", x"7876", x"7875", x"7874", 
    x"7873", x"7872", x"7870", x"786f", x"786e", x"786d", x"786c", x"786b", 
    x"786a", x"7869", x"7868", x"7867", x"7866", x"7865", x"7864", x"7863", 
    x"7862", x"7860", x"785f", x"785e", x"785d", x"785c", x"785b", x"785a", 
    x"7859", x"7858", x"7857", x"7856", x"7855", x"7854", x"7853", x"7852", 
    x"7850", x"784f", x"784e", x"784d", x"784c", x"784b", x"784a", x"7849", 
    x"7848", x"7847", x"7846", x"7845", x"7844", x"7842", x"7841", x"7840", 
    x"783f", x"783e", x"783d", x"783c", x"783b", x"783a", x"7839", x"7838", 
    x"7837", x"7836", x"7834", x"7833", x"7832", x"7831", x"7830", x"782f", 
    x"782e", x"782d", x"782c", x"782b", x"782a", x"7829", x"7828", x"7826", 
    x"7825", x"7824", x"7823", x"7822", x"7821", x"7820", x"781f", x"781e", 
    x"781d", x"781c", x"781a", x"7819", x"7818", x"7817", x"7816", x"7815", 
    x"7814", x"7813", x"7812", x"7811", x"7810", x"780f", x"780d", x"780c", 
    x"780b", x"780a", x"7809", x"7808", x"7807", x"7806", x"7805", x"7804", 
    x"7803", x"7801", x"7800", x"77ff", x"77fe", x"77fd", x"77fc", x"77fb", 
    x"77fa", x"77f9", x"77f8", x"77f7", x"77f5", x"77f4", x"77f3", x"77f2", 
    x"77f1", x"77f0", x"77ef", x"77ee", x"77ed", x"77ec", x"77ea", x"77e9", 
    x"77e8", x"77e7", x"77e6", x"77e5", x"77e4", x"77e3", x"77e2", x"77e1", 
    x"77df", x"77de", x"77dd", x"77dc", x"77db", x"77da", x"77d9", x"77d8", 
    x"77d7", x"77d6", x"77d4", x"77d3", x"77d2", x"77d1", x"77d0", x"77cf", 
    x"77ce", x"77cd", x"77cc", x"77ca", x"77c9", x"77c8", x"77c7", x"77c6", 
    x"77c5", x"77c4", x"77c3", x"77c2", x"77c0", x"77bf", x"77be", x"77bd", 
    x"77bc", x"77bb", x"77ba", x"77b9", x"77b8", x"77b6", x"77b5", x"77b4", 
    x"77b3", x"77b2", x"77b1", x"77b0", x"77af", x"77ae", x"77ac", x"77ab", 
    x"77aa", x"77a9", x"77a8", x"77a7", x"77a6", x"77a5", x"77a4", x"77a2", 
    x"77a1", x"77a0", x"779f", x"779e", x"779d", x"779c", x"779b", x"7799", 
    x"7798", x"7797", x"7796", x"7795", x"7794", x"7793", x"7792", x"7791", 
    x"778f", x"778e", x"778d", x"778c", x"778b", x"778a", x"7789", x"7788", 
    x"7786", x"7785", x"7784", x"7783", x"7782", x"7781", x"7780", x"777f", 
    x"777d", x"777c", x"777b", x"777a", x"7779", x"7778", x"7777", x"7776", 
    x"7774", x"7773", x"7772", x"7771", x"7770", x"776f", x"776e", x"776d", 
    x"776b", x"776a", x"7769", x"7768", x"7767", x"7766", x"7765", x"7763", 
    x"7762", x"7761", x"7760", x"775f", x"775e", x"775d", x"775c", x"775a", 
    x"7759", x"7758", x"7757", x"7756", x"7755", x"7754", x"7752", x"7751", 
    x"7750", x"774f", x"774e", x"774d", x"774c", x"774a", x"7749", x"7748", 
    x"7747", x"7746", x"7745", x"7744", x"7742", x"7741", x"7740", x"773f", 
    x"773e", x"773d", x"773c", x"773a", x"7739", x"7738", x"7737", x"7736", 
    x"7735", x"7734", x"7732", x"7731", x"7730", x"772f", x"772e", x"772d", 
    x"772c", x"772a", x"7729", x"7728", x"7727", x"7726", x"7725", x"7724", 
    x"7722", x"7721", x"7720", x"771f", x"771e", x"771d", x"771c", x"771a", 
    x"7719", x"7718", x"7717", x"7716", x"7715", x"7713", x"7712", x"7711", 
    x"7710", x"770f", x"770e", x"770d", x"770b", x"770a", x"7709", x"7708", 
    x"7707", x"7706", x"7704", x"7703", x"7702", x"7701", x"7700", x"76ff", 
    x"76fe", x"76fc", x"76fb", x"76fa", x"76f9", x"76f8", x"76f7", x"76f5", 
    x"76f4", x"76f3", x"76f2", x"76f1", x"76f0", x"76ee", x"76ed", x"76ec", 
    x"76eb", x"76ea", x"76e9", x"76e7", x"76e6", x"76e5", x"76e4", x"76e3", 
    x"76e2", x"76e1", x"76df", x"76de", x"76dd", x"76dc", x"76db", x"76da", 
    x"76d8", x"76d7", x"76d6", x"76d5", x"76d4", x"76d3", x"76d1", x"76d0", 
    x"76cf", x"76ce", x"76cd", x"76cc", x"76ca", x"76c9", x"76c8", x"76c7", 
    x"76c6", x"76c4", x"76c3", x"76c2", x"76c1", x"76c0", x"76bf", x"76bd", 
    x"76bc", x"76bb", x"76ba", x"76b9", x"76b8", x"76b6", x"76b5", x"76b4", 
    x"76b3", x"76b2", x"76b1", x"76af", x"76ae", x"76ad", x"76ac", x"76ab", 
    x"76a9", x"76a8", x"76a7", x"76a6", x"76a5", x"76a4", x"76a2", x"76a1", 
    x"76a0", x"769f", x"769e", x"769d", x"769b", x"769a", x"7699", x"7698", 
    x"7697", x"7695", x"7694", x"7693", x"7692", x"7691", x"768f", x"768e", 
    x"768d", x"768c", x"768b", x"768a", x"7688", x"7687", x"7686", x"7685", 
    x"7684", x"7682", x"7681", x"7680", x"767f", x"767e", x"767d", x"767b", 
    x"767a", x"7679", x"7678", x"7677", x"7675", x"7674", x"7673", x"7672", 
    x"7671", x"766f", x"766e", x"766d", x"766c", x"766b", x"7669", x"7668", 
    x"7667", x"7666", x"7665", x"7664", x"7662", x"7661", x"7660", x"765f", 
    x"765e", x"765c", x"765b", x"765a", x"7659", x"7658", x"7656", x"7655", 
    x"7654", x"7653", x"7652", x"7650", x"764f", x"764e", x"764d", x"764c", 
    x"764a", x"7649", x"7648", x"7647", x"7646", x"7644", x"7643", x"7642", 
    x"7641", x"7640", x"763e", x"763d", x"763c", x"763b", x"763a", x"7638", 
    x"7637", x"7636", x"7635", x"7634", x"7632", x"7631", x"7630", x"762f", 
    x"762d", x"762c", x"762b", x"762a", x"7629", x"7627", x"7626", x"7625", 
    x"7624", x"7623", x"7621", x"7620", x"761f", x"761e", x"761d", x"761b", 
    x"761a", x"7619", x"7618", x"7617", x"7615", x"7614", x"7613", x"7612", 
    x"7610", x"760f", x"760e", x"760d", x"760c", x"760a", x"7609", x"7608", 
    x"7607", x"7606", x"7604", x"7603", x"7602", x"7601", x"75ff", x"75fe", 
    x"75fd", x"75fc", x"75fb", x"75f9", x"75f8", x"75f7", x"75f6", x"75f4", 
    x"75f3", x"75f2", x"75f1", x"75f0", x"75ee", x"75ed", x"75ec", x"75eb", 
    x"75e9", x"75e8", x"75e7", x"75e6", x"75e5", x"75e3", x"75e2", x"75e1", 
    x"75e0", x"75de", x"75dd", x"75dc", x"75db", x"75da", x"75d8", x"75d7", 
    x"75d6", x"75d5", x"75d3", x"75d2", x"75d1", x"75d0", x"75cf", x"75cd", 
    x"75cc", x"75cb", x"75ca", x"75c8", x"75c7", x"75c6", x"75c5", x"75c3", 
    x"75c2", x"75c1", x"75c0", x"75bf", x"75bd", x"75bc", x"75bb", x"75ba", 
    x"75b8", x"75b7", x"75b6", x"75b5", x"75b3", x"75b2", x"75b1", x"75b0", 
    x"75ae", x"75ad", x"75ac", x"75ab", x"75aa", x"75a8", x"75a7", x"75a6", 
    x"75a5", x"75a3", x"75a2", x"75a1", x"75a0", x"759e", x"759d", x"759c", 
    x"759b", x"7599", x"7598", x"7597", x"7596", x"7594", x"7593", x"7592", 
    x"7591", x"7590", x"758e", x"758d", x"758c", x"758b", x"7589", x"7588", 
    x"7587", x"7586", x"7584", x"7583", x"7582", x"7581", x"757f", x"757e", 
    x"757d", x"757c", x"757a", x"7579", x"7578", x"7577", x"7575", x"7574", 
    x"7573", x"7572", x"7570", x"756f", x"756e", x"756d", x"756b", x"756a", 
    x"7569", x"7568", x"7566", x"7565", x"7564", x"7563", x"7561", x"7560", 
    x"755f", x"755e", x"755c", x"755b", x"755a", x"7559", x"7557", x"7556", 
    x"7555", x"7554", x"7552", x"7551", x"7550", x"754f", x"754d", x"754c", 
    x"754b", x"754a", x"7548", x"7547", x"7546", x"7544", x"7543", x"7542", 
    x"7541", x"753f", x"753e", x"753d", x"753c", x"753a", x"7539", x"7538", 
    x"7537", x"7535", x"7534", x"7533", x"7532", x"7530", x"752f", x"752e", 
    x"752d", x"752b", x"752a", x"7529", x"7527", x"7526", x"7525", x"7524", 
    x"7522", x"7521", x"7520", x"751f", x"751d", x"751c", x"751b", x"751a", 
    x"7518", x"7517", x"7516", x"7514", x"7513", x"7512", x"7511", x"750f", 
    x"750e", x"750d", x"750c", x"750a", x"7509", x"7508", x"7506", x"7505", 
    x"7504", x"7503", x"7501", x"7500", x"74ff", x"74fe", x"74fc", x"74fb", 
    x"74fa", x"74f8", x"74f7", x"74f6", x"74f5", x"74f3", x"74f2", x"74f1", 
    x"74f0", x"74ee", x"74ed", x"74ec", x"74ea", x"74e9", x"74e8", x"74e7", 
    x"74e5", x"74e4", x"74e3", x"74e1", x"74e0", x"74df", x"74de", x"74dc", 
    x"74db", x"74da", x"74d8", x"74d7", x"74d6", x"74d5", x"74d3", x"74d2", 
    x"74d1", x"74cf", x"74ce", x"74cd", x"74cc", x"74ca", x"74c9", x"74c8", 
    x"74c6", x"74c5", x"74c4", x"74c3", x"74c1", x"74c0", x"74bf", x"74bd", 
    x"74bc", x"74bb", x"74ba", x"74b8", x"74b7", x"74b6", x"74b4", x"74b3", 
    x"74b2", x"74b1", x"74af", x"74ae", x"74ad", x"74ab", x"74aa", x"74a9", 
    x"74a8", x"74a6", x"74a5", x"74a4", x"74a2", x"74a1", x"74a0", x"749e", 
    x"749d", x"749c", x"749b", x"7499", x"7498", x"7497", x"7495", x"7494", 
    x"7493", x"7492", x"7490", x"748f", x"748e", x"748c", x"748b", x"748a", 
    x"7488", x"7487", x"7486", x"7485", x"7483", x"7482", x"7481", x"747f", 
    x"747e", x"747d", x"747b", x"747a", x"7479", x"7478", x"7476", x"7475", 
    x"7474", x"7472", x"7471", x"7470", x"746e", x"746d", x"746c", x"746a", 
    x"7469", x"7468", x"7467", x"7465", x"7464", x"7463", x"7461", x"7460", 
    x"745f", x"745d", x"745c", x"745b", x"7459", x"7458", x"7457", x"7456", 
    x"7454", x"7453", x"7452", x"7450", x"744f", x"744e", x"744c", x"744b", 
    x"744a", x"7448", x"7447", x"7446", x"7444", x"7443", x"7442", x"7441", 
    x"743f", x"743e", x"743d", x"743b", x"743a", x"7439", x"7437", x"7436", 
    x"7435", x"7433", x"7432", x"7431", x"742f", x"742e", x"742d", x"742b", 
    x"742a", x"7429", x"7428", x"7426", x"7425", x"7424", x"7422", x"7421", 
    x"7420", x"741e", x"741d", x"741c", x"741a", x"7419", x"7418", x"7416", 
    x"7415", x"7414", x"7412", x"7411", x"7410", x"740e", x"740d", x"740c", 
    x"740a", x"7409", x"7408", x"7406", x"7405", x"7404", x"7402", x"7401", 
    x"7400", x"73fe", x"73fd", x"73fc", x"73fa", x"73f9", x"73f8", x"73f7", 
    x"73f5", x"73f4", x"73f3", x"73f1", x"73f0", x"73ef", x"73ed", x"73ec", 
    x"73eb", x"73e9", x"73e8", x"73e7", x"73e5", x"73e4", x"73e3", x"73e1", 
    x"73e0", x"73df", x"73dd", x"73dc", x"73db", x"73d9", x"73d8", x"73d7", 
    x"73d5", x"73d4", x"73d3", x"73d1", x"73d0", x"73ce", x"73cd", x"73cc", 
    x"73ca", x"73c9", x"73c8", x"73c6", x"73c5", x"73c4", x"73c2", x"73c1", 
    x"73c0", x"73be", x"73bd", x"73bc", x"73ba", x"73b9", x"73b8", x"73b6", 
    x"73b5", x"73b4", x"73b2", x"73b1", x"73b0", x"73ae", x"73ad", x"73ac", 
    x"73aa", x"73a9", x"73a8", x"73a6", x"73a5", x"73a4", x"73a2", x"73a1", 
    x"739f", x"739e", x"739d", x"739b", x"739a", x"7399", x"7397", x"7396", 
    x"7395", x"7393", x"7392", x"7391", x"738f", x"738e", x"738d", x"738b", 
    x"738a", x"7389", x"7387", x"7386", x"7384", x"7383", x"7382", x"7380", 
    x"737f", x"737e", x"737c", x"737b", x"737a", x"7378", x"7377", x"7376", 
    x"7374", x"7373", x"7372", x"7370", x"736f", x"736d", x"736c", x"736b", 
    x"7369", x"7368", x"7367", x"7365", x"7364", x"7363", x"7361", x"7360", 
    x"735e", x"735d", x"735c", x"735a", x"7359", x"7358", x"7356", x"7355", 
    x"7354", x"7352", x"7351", x"7350", x"734e", x"734d", x"734b", x"734a", 
    x"7349", x"7347", x"7346", x"7345", x"7343", x"7342", x"7340", x"733f", 
    x"733e", x"733c", x"733b", x"733a", x"7338", x"7337", x"7336", x"7334", 
    x"7333", x"7331", x"7330", x"732f", x"732d", x"732c", x"732b", x"7329", 
    x"7328", x"7326", x"7325", x"7324", x"7322", x"7321", x"7320", x"731e", 
    x"731d", x"731c", x"731a", x"7319", x"7317", x"7316", x"7315", x"7313", 
    x"7312", x"7311", x"730f", x"730e", x"730c", x"730b", x"730a", x"7308", 
    x"7307", x"7305", x"7304", x"7303", x"7301", x"7300", x"72ff", x"72fd", 
    x"72fc", x"72fa", x"72f9", x"72f8", x"72f6", x"72f5", x"72f4", x"72f2", 
    x"72f1", x"72ef", x"72ee", x"72ed", x"72eb", x"72ea", x"72e8", x"72e7", 
    x"72e6", x"72e4", x"72e3", x"72e2", x"72e0", x"72df", x"72dd", x"72dc", 
    x"72db", x"72d9", x"72d8", x"72d6", x"72d5", x"72d4", x"72d2", x"72d1", 
    x"72d0", x"72ce", x"72cd", x"72cb", x"72ca", x"72c9", x"72c7", x"72c6", 
    x"72c4", x"72c3", x"72c2", x"72c0", x"72bf", x"72bd", x"72bc", x"72bb", 
    x"72b9", x"72b8", x"72b6", x"72b5", x"72b4", x"72b2", x"72b1", x"72b0", 
    x"72ae", x"72ad", x"72ab", x"72aa", x"72a9", x"72a7", x"72a6", x"72a4", 
    x"72a3", x"72a2", x"72a0", x"729f", x"729d", x"729c", x"729b", x"7299", 
    x"7298", x"7296", x"7295", x"7294", x"7292", x"7291", x"728f", x"728e", 
    x"728d", x"728b", x"728a", x"7288", x"7287", x"7286", x"7284", x"7283", 
    x"7281", x"7280", x"727f", x"727d", x"727c", x"727a", x"7279", x"7278", 
    x"7276", x"7275", x"7273", x"7272", x"7270", x"726f", x"726e", x"726c", 
    x"726b", x"7269", x"7268", x"7267", x"7265", x"7264", x"7262", x"7261", 
    x"7260", x"725e", x"725d", x"725b", x"725a", x"7259", x"7257", x"7256", 
    x"7254", x"7253", x"7251", x"7250", x"724f", x"724d", x"724c", x"724a", 
    x"7249", x"7248", x"7246", x"7245", x"7243", x"7242", x"7240", x"723f", 
    x"723e", x"723c", x"723b", x"7239", x"7238", x"7237", x"7235", x"7234", 
    x"7232", x"7231", x"722f", x"722e", x"722d", x"722b", x"722a", x"7228", 
    x"7227", x"7226", x"7224", x"7223", x"7221", x"7220", x"721e", x"721d", 
    x"721c", x"721a", x"7219", x"7217", x"7216", x"7214", x"7213", x"7212", 
    x"7210", x"720f", x"720d", x"720c", x"720a", x"7209", x"7208", x"7206", 
    x"7205", x"7203", x"7202", x"7200", x"71ff", x"71fe", x"71fc", x"71fb", 
    x"71f9", x"71f8", x"71f6", x"71f5", x"71f4", x"71f2", x"71f1", x"71ef", 
    x"71ee", x"71ec", x"71eb", x"71ea", x"71e8", x"71e7", x"71e5", x"71e4", 
    x"71e2", x"71e1", x"71e0", x"71de", x"71dd", x"71db", x"71da", x"71d8", 
    x"71d7", x"71d6", x"71d4", x"71d3", x"71d1", x"71d0", x"71ce", x"71cd", 
    x"71cb", x"71ca", x"71c9", x"71c7", x"71c6", x"71c4", x"71c3", x"71c1", 
    x"71c0", x"71be", x"71bd", x"71bc", x"71ba", x"71b9", x"71b7", x"71b6", 
    x"71b4", x"71b3", x"71b2", x"71b0", x"71af", x"71ad", x"71ac", x"71aa", 
    x"71a9", x"71a7", x"71a6", x"71a5", x"71a3", x"71a2", x"71a0", x"719f", 
    x"719d", x"719c", x"719a", x"7199", x"7197", x"7196", x"7195", x"7193", 
    x"7192", x"7190", x"718f", x"718d", x"718c", x"718a", x"7189", x"7188", 
    x"7186", x"7185", x"7183", x"7182", x"7180", x"717f", x"717d", x"717c", 
    x"717a", x"7179", x"7178", x"7176", x"7175", x"7173", x"7172", x"7170", 
    x"716f", x"716d", x"716c", x"716a", x"7169", x"7168", x"7166", x"7165", 
    x"7163", x"7162", x"7160", x"715f", x"715d", x"715c", x"715a", x"7159", 
    x"7158", x"7156", x"7155", x"7153", x"7152", x"7150", x"714f", x"714d", 
    x"714c", x"714a", x"7149", x"7147", x"7146", x"7145", x"7143", x"7142", 
    x"7140", x"713f", x"713d", x"713c", x"713a", x"7139", x"7137", x"7136", 
    x"7134", x"7133", x"7131", x"7130", x"712f", x"712d", x"712c", x"712a", 
    x"7129", x"7127", x"7126", x"7124", x"7123", x"7121", x"7120", x"711e", 
    x"711d", x"711b", x"711a", x"7119", x"7117", x"7116", x"7114", x"7113", 
    x"7111", x"7110", x"710e", x"710d", x"710b", x"710a", x"7108", x"7107", 
    x"7105", x"7104", x"7102", x"7101", x"70ff", x"70fe", x"70fd", x"70fb", 
    x"70fa", x"70f8", x"70f7", x"70f5", x"70f4", x"70f2", x"70f1", x"70ef", 
    x"70ee", x"70ec", x"70eb", x"70e9", x"70e8", x"70e6", x"70e5", x"70e3", 
    x"70e2", x"70e0", x"70df", x"70dd", x"70dc", x"70db", x"70d9", x"70d8", 
    x"70d6", x"70d5", x"70d3", x"70d2", x"70d0", x"70cf", x"70cd", x"70cc", 
    x"70ca", x"70c9", x"70c7", x"70c6", x"70c4", x"70c3", x"70c1", x"70c0", 
    x"70be", x"70bd", x"70bb", x"70ba", x"70b8", x"70b7", x"70b5", x"70b4", 
    x"70b2", x"70b1", x"70af", x"70ae", x"70ac", x"70ab", x"70a9", x"70a8", 
    x"70a6", x"70a5", x"70a3", x"70a2", x"70a0", x"709f", x"709e", x"709c", 
    x"709b", x"7099", x"7098", x"7096", x"7095", x"7093", x"7092", x"7090", 
    x"708f", x"708d", x"708c", x"708a", x"7089", x"7087", x"7086", x"7084", 
    x"7083", x"7081", x"7080", x"707e", x"707d", x"707b", x"707a", x"7078", 
    x"7077", x"7075", x"7074", x"7072", x"7071", x"706f", x"706e", x"706c", 
    x"706b", x"7069", x"7068", x"7066", x"7065", x"7063", x"7062", x"7060", 
    x"705f", x"705d", x"705c", x"705a", x"7059", x"7057", x"7056", x"7054", 
    x"7053", x"7051", x"7050", x"704e", x"704c", x"704b", x"7049", x"7048", 
    x"7046", x"7045", x"7043", x"7042", x"7040", x"703f", x"703d", x"703c", 
    x"703a", x"7039", x"7037", x"7036", x"7034", x"7033", x"7031", x"7030", 
    x"702e", x"702d", x"702b", x"702a", x"7028", x"7027", x"7025", x"7024", 
    x"7022", x"7021", x"701f", x"701e", x"701c", x"701b", x"7019", x"7018", 
    x"7016", x"7015", x"7013", x"7012", x"7010", x"700e", x"700d", x"700b", 
    x"700a", x"7008", x"7007", x"7005", x"7004", x"7002", x"7001", x"6fff", 
    x"6ffe", x"6ffc", x"6ffb", x"6ff9", x"6ff8", x"6ff6", x"6ff5", x"6ff3", 
    x"6ff2", x"6ff0", x"6fef", x"6fed", x"6feb", x"6fea", x"6fe8", x"6fe7", 
    x"6fe5", x"6fe4", x"6fe2", x"6fe1", x"6fdf", x"6fde", x"6fdc", x"6fdb", 
    x"6fd9", x"6fd8", x"6fd6", x"6fd5", x"6fd3", x"6fd2", x"6fd0", x"6fce", 
    x"6fcd", x"6fcb", x"6fca", x"6fc8", x"6fc7", x"6fc5", x"6fc4", x"6fc2", 
    x"6fc1", x"6fbf", x"6fbe", x"6fbc", x"6fbb", x"6fb9", x"6fb8", x"6fb6", 
    x"6fb4", x"6fb3", x"6fb1", x"6fb0", x"6fae", x"6fad", x"6fab", x"6faa", 
    x"6fa8", x"6fa7", x"6fa5", x"6fa4", x"6fa2", x"6fa0", x"6f9f", x"6f9d", 
    x"6f9c", x"6f9a", x"6f99", x"6f97", x"6f96", x"6f94", x"6f93", x"6f91", 
    x"6f90", x"6f8e", x"6f8c", x"6f8b", x"6f89", x"6f88", x"6f86", x"6f85", 
    x"6f83", x"6f82", x"6f80", x"6f7f", x"6f7d", x"6f7c", x"6f7a", x"6f78", 
    x"6f77", x"6f75", x"6f74", x"6f72", x"6f71", x"6f6f", x"6f6e", x"6f6c", 
    x"6f6b", x"6f69", x"6f67", x"6f66", x"6f64", x"6f63", x"6f61", x"6f60", 
    x"6f5e", x"6f5d", x"6f5b", x"6f59", x"6f58", x"6f56", x"6f55", x"6f53", 
    x"6f52", x"6f50", x"6f4f", x"6f4d", x"6f4c", x"6f4a", x"6f48", x"6f47", 
    x"6f45", x"6f44", x"6f42", x"6f41", x"6f3f", x"6f3e", x"6f3c", x"6f3a", 
    x"6f39", x"6f37", x"6f36", x"6f34", x"6f33", x"6f31", x"6f30", x"6f2e", 
    x"6f2c", x"6f2b", x"6f29", x"6f28", x"6f26", x"6f25", x"6f23", x"6f22", 
    x"6f20", x"6f1e", x"6f1d", x"6f1b", x"6f1a", x"6f18", x"6f17", x"6f15", 
    x"6f14", x"6f12", x"6f10", x"6f0f", x"6f0d", x"6f0c", x"6f0a", x"6f09", 
    x"6f07", x"6f05", x"6f04", x"6f02", x"6f01", x"6eff", x"6efe", x"6efc", 
    x"6efb", x"6ef9", x"6ef7", x"6ef6", x"6ef4", x"6ef3", x"6ef1", x"6ef0", 
    x"6eee", x"6eec", x"6eeb", x"6ee9", x"6ee8", x"6ee6", x"6ee5", x"6ee3", 
    x"6ee1", x"6ee0", x"6ede", x"6edd", x"6edb", x"6eda", x"6ed8", x"6ed6", 
    x"6ed5", x"6ed3", x"6ed2", x"6ed0", x"6ecf", x"6ecd", x"6ecb", x"6eca", 
    x"6ec8", x"6ec7", x"6ec5", x"6ec4", x"6ec2", x"6ec0", x"6ebf", x"6ebd", 
    x"6ebc", x"6eba", x"6eb9", x"6eb7", x"6eb5", x"6eb4", x"6eb2", x"6eb1", 
    x"6eaf", x"6ead", x"6eac", x"6eaa", x"6ea9", x"6ea7", x"6ea6", x"6ea4", 
    x"6ea2", x"6ea1", x"6e9f", x"6e9e", x"6e9c", x"6e9b", x"6e99", x"6e97", 
    x"6e96", x"6e94", x"6e93", x"6e91", x"6e8f", x"6e8e", x"6e8c", x"6e8b", 
    x"6e89", x"6e88", x"6e86", x"6e84", x"6e83", x"6e81", x"6e80", x"6e7e", 
    x"6e7c", x"6e7b", x"6e79", x"6e78", x"6e76", x"6e75", x"6e73", x"6e71", 
    x"6e70", x"6e6e", x"6e6d", x"6e6b", x"6e69", x"6e68", x"6e66", x"6e65", 
    x"6e63", x"6e61", x"6e60", x"6e5e", x"6e5d", x"6e5b", x"6e59", x"6e58", 
    x"6e56", x"6e55", x"6e53", x"6e52", x"6e50", x"6e4e", x"6e4d", x"6e4b", 
    x"6e4a", x"6e48", x"6e46", x"6e45", x"6e43", x"6e42", x"6e40", x"6e3e", 
    x"6e3d", x"6e3b", x"6e3a", x"6e38", x"6e36", x"6e35", x"6e33", x"6e32", 
    x"6e30", x"6e2e", x"6e2d", x"6e2b", x"6e2a", x"6e28", x"6e26", x"6e25", 
    x"6e23", x"6e22", x"6e20", x"6e1e", x"6e1d", x"6e1b", x"6e1a", x"6e18", 
    x"6e16", x"6e15", x"6e13", x"6e12", x"6e10", x"6e0e", x"6e0d", x"6e0b", 
    x"6e0a", x"6e08", x"6e06", x"6e05", x"6e03", x"6e02", x"6e00", x"6dfe", 
    x"6dfd", x"6dfb", x"6dfa", x"6df8", x"6df6", x"6df5", x"6df3", x"6df1", 
    x"6df0", x"6dee", x"6ded", x"6deb", x"6de9", x"6de8", x"6de6", x"6de5", 
    x"6de3", x"6de1", x"6de0", x"6dde", x"6ddd", x"6ddb", x"6dd9", x"6dd8", 
    x"6dd6", x"6dd4", x"6dd3", x"6dd1", x"6dd0", x"6dce", x"6dcc", x"6dcb", 
    x"6dc9", x"6dc8", x"6dc6", x"6dc4", x"6dc3", x"6dc1", x"6dbf", x"6dbe", 
    x"6dbc", x"6dbb", x"6db9", x"6db7", x"6db6", x"6db4", x"6db3", x"6db1", 
    x"6daf", x"6dae", x"6dac", x"6daa", x"6da9", x"6da7", x"6da6", x"6da4", 
    x"6da2", x"6da1", x"6d9f", x"6d9d", x"6d9c", x"6d9a", x"6d99", x"6d97", 
    x"6d95", x"6d94", x"6d92", x"6d91", x"6d8f", x"6d8d", x"6d8c", x"6d8a", 
    x"6d88", x"6d87", x"6d85", x"6d84", x"6d82", x"6d80", x"6d7f", x"6d7d", 
    x"6d7b", x"6d7a", x"6d78", x"6d76", x"6d75", x"6d73", x"6d72", x"6d70", 
    x"6d6e", x"6d6d", x"6d6b", x"6d69", x"6d68", x"6d66", x"6d65", x"6d63", 
    x"6d61", x"6d60", x"6d5e", x"6d5c", x"6d5b", x"6d59", x"6d58", x"6d56", 
    x"6d54", x"6d53", x"6d51", x"6d4f", x"6d4e", x"6d4c", x"6d4a", x"6d49", 
    x"6d47", x"6d46", x"6d44", x"6d42", x"6d41", x"6d3f", x"6d3d", x"6d3c", 
    x"6d3a", x"6d38", x"6d37", x"6d35", x"6d34", x"6d32", x"6d30", x"6d2f", 
    x"6d2d", x"6d2b", x"6d2a", x"6d28", x"6d26", x"6d25", x"6d23", x"6d21", 
    x"6d20", x"6d1e", x"6d1d", x"6d1b", x"6d19", x"6d18", x"6d16", x"6d14", 
    x"6d13", x"6d11", x"6d0f", x"6d0e", x"6d0c", x"6d0a", x"6d09", x"6d07", 
    x"6d06", x"6d04", x"6d02", x"6d01", x"6cff", x"6cfd", x"6cfc", x"6cfa", 
    x"6cf8", x"6cf7", x"6cf5", x"6cf3", x"6cf2", x"6cf0", x"6cee", x"6ced", 
    x"6ceb", x"6cea", x"6ce8", x"6ce6", x"6ce5", x"6ce3", x"6ce1", x"6ce0", 
    x"6cde", x"6cdc", x"6cdb", x"6cd9", x"6cd7", x"6cd6", x"6cd4", x"6cd2", 
    x"6cd1", x"6ccf", x"6ccd", x"6ccc", x"6cca", x"6cc8", x"6cc7", x"6cc5", 
    x"6cc3", x"6cc2", x"6cc0", x"6cbf", x"6cbd", x"6cbb", x"6cba", x"6cb8", 
    x"6cb6", x"6cb5", x"6cb3", x"6cb1", x"6cb0", x"6cae", x"6cac", x"6cab", 
    x"6ca9", x"6ca7", x"6ca6", x"6ca4", x"6ca2", x"6ca1", x"6c9f", x"6c9d", 
    x"6c9c", x"6c9a", x"6c98", x"6c97", x"6c95", x"6c93", x"6c92", x"6c90", 
    x"6c8e", x"6c8d", x"6c8b", x"6c89", x"6c88", x"6c86", x"6c84", x"6c83", 
    x"6c81", x"6c7f", x"6c7e", x"6c7c", x"6c7a", x"6c79", x"6c77", x"6c75", 
    x"6c74", x"6c72", x"6c70", x"6c6f", x"6c6d", x"6c6b", x"6c6a", x"6c68", 
    x"6c66", x"6c65", x"6c63", x"6c61", x"6c60", x"6c5e", x"6c5c", x"6c5b", 
    x"6c59", x"6c57", x"6c56", x"6c54", x"6c52", x"6c51", x"6c4f", x"6c4d", 
    x"6c4c", x"6c4a", x"6c48", x"6c47", x"6c45", x"6c43", x"6c42", x"6c40", 
    x"6c3e", x"6c3c", x"6c3b", x"6c39", x"6c37", x"6c36", x"6c34", x"6c32", 
    x"6c31", x"6c2f", x"6c2d", x"6c2c", x"6c2a", x"6c28", x"6c27", x"6c25", 
    x"6c23", x"6c22", x"6c20", x"6c1e", x"6c1d", x"6c1b", x"6c19", x"6c18", 
    x"6c16", x"6c14", x"6c12", x"6c11", x"6c0f", x"6c0d", x"6c0c", x"6c0a", 
    x"6c08", x"6c07", x"6c05", x"6c03", x"6c02", x"6c00", x"6bfe", x"6bfd", 
    x"6bfb", x"6bf9", x"6bf8", x"6bf6", x"6bf4", x"6bf2", x"6bf1", x"6bef", 
    x"6bed", x"6bec", x"6bea", x"6be8", x"6be7", x"6be5", x"6be3", x"6be2", 
    x"6be0", x"6bde", x"6bdd", x"6bdb", x"6bd9", x"6bd7", x"6bd6", x"6bd4", 
    x"6bd2", x"6bd1", x"6bcf", x"6bcd", x"6bcc", x"6bca", x"6bc8", x"6bc6", 
    x"6bc5", x"6bc3", x"6bc1", x"6bc0", x"6bbe", x"6bbc", x"6bbb", x"6bb9", 
    x"6bb7", x"6bb6", x"6bb4", x"6bb2", x"6bb0", x"6baf", x"6bad", x"6bab", 
    x"6baa", x"6ba8", x"6ba6", x"6ba5", x"6ba3", x"6ba1", x"6b9f", x"6b9e", 
    x"6b9c", x"6b9a", x"6b99", x"6b97", x"6b95", x"6b94", x"6b92", x"6b90", 
    x"6b8e", x"6b8d", x"6b8b", x"6b89", x"6b88", x"6b86", x"6b84", x"6b83", 
    x"6b81", x"6b7f", x"6b7d", x"6b7c", x"6b7a", x"6b78", x"6b77", x"6b75", 
    x"6b73", x"6b71", x"6b70", x"6b6e", x"6b6c", x"6b6b", x"6b69", x"6b67", 
    x"6b65", x"6b64", x"6b62", x"6b60", x"6b5f", x"6b5d", x"6b5b", x"6b5a", 
    x"6b58", x"6b56", x"6b54", x"6b53", x"6b51", x"6b4f", x"6b4e", x"6b4c", 
    x"6b4a", x"6b48", x"6b47", x"6b45", x"6b43", x"6b42", x"6b40", x"6b3e", 
    x"6b3c", x"6b3b", x"6b39", x"6b37", x"6b36", x"6b34", x"6b32", x"6b30", 
    x"6b2f", x"6b2d", x"6b2b", x"6b2a", x"6b28", x"6b26", x"6b24", x"6b23", 
    x"6b21", x"6b1f", x"6b1d", x"6b1c", x"6b1a", x"6b18", x"6b17", x"6b15", 
    x"6b13", x"6b11", x"6b10", x"6b0e", x"6b0c", x"6b0b", x"6b09", x"6b07", 
    x"6b05", x"6b04", x"6b02", x"6b00", x"6afe", x"6afd", x"6afb", x"6af9", 
    x"6af8", x"6af6", x"6af4", x"6af2", x"6af1", x"6aef", x"6aed", x"6aec", 
    x"6aea", x"6ae8", x"6ae6", x"6ae5", x"6ae3", x"6ae1", x"6adf", x"6ade", 
    x"6adc", x"6ada", x"6ad8", x"6ad7", x"6ad5", x"6ad3", x"6ad2", x"6ad0", 
    x"6ace", x"6acc", x"6acb", x"6ac9", x"6ac7", x"6ac5", x"6ac4", x"6ac2", 
    x"6ac0", x"6abf", x"6abd", x"6abb", x"6ab9", x"6ab8", x"6ab6", x"6ab4", 
    x"6ab2", x"6ab1", x"6aaf", x"6aad", x"6aab", x"6aaa", x"6aa8", x"6aa6", 
    x"6aa4", x"6aa3", x"6aa1", x"6a9f", x"6a9e", x"6a9c", x"6a9a", x"6a98", 
    x"6a97", x"6a95", x"6a93", x"6a91", x"6a90", x"6a8e", x"6a8c", x"6a8a", 
    x"6a89", x"6a87", x"6a85", x"6a83", x"6a82", x"6a80", x"6a7e", x"6a7c", 
    x"6a7b", x"6a79", x"6a77", x"6a75", x"6a74", x"6a72", x"6a70", x"6a6f", 
    x"6a6d", x"6a6b", x"6a69", x"6a68", x"6a66", x"6a64", x"6a62", x"6a61", 
    x"6a5f", x"6a5d", x"6a5b", x"6a5a", x"6a58", x"6a56", x"6a54", x"6a53", 
    x"6a51", x"6a4f", x"6a4d", x"6a4c", x"6a4a", x"6a48", x"6a46", x"6a45", 
    x"6a43", x"6a41", x"6a3f", x"6a3e", x"6a3c", x"6a3a", x"6a38", x"6a37", 
    x"6a35", x"6a33", x"6a31", x"6a30", x"6a2e", x"6a2c", x"6a2a", x"6a29", 
    x"6a27", x"6a25", x"6a23", x"6a21", x"6a20", x"6a1e", x"6a1c", x"6a1a", 
    x"6a19", x"6a17", x"6a15", x"6a13", x"6a12", x"6a10", x"6a0e", x"6a0c", 
    x"6a0b", x"6a09", x"6a07", x"6a05", x"6a04", x"6a02", x"6a00", x"69fe", 
    x"69fd", x"69fb", x"69f9", x"69f7", x"69f6", x"69f4", x"69f2", x"69f0", 
    x"69ee", x"69ed", x"69eb", x"69e9", x"69e7", x"69e6", x"69e4", x"69e2", 
    x"69e0", x"69df", x"69dd", x"69db", x"69d9", x"69d8", x"69d6", x"69d4", 
    x"69d2", x"69d0", x"69cf", x"69cd", x"69cb", x"69c9", x"69c8", x"69c6", 
    x"69c4", x"69c2", x"69c1", x"69bf", x"69bd", x"69bb", x"69b9", x"69b8", 
    x"69b6", x"69b4", x"69b2", x"69b1", x"69af", x"69ad", x"69ab", x"69a9", 
    x"69a8", x"69a6", x"69a4", x"69a2", x"69a1", x"699f", x"699d", x"699b", 
    x"699a", x"6998", x"6996", x"6994", x"6992", x"6991", x"698f", x"698d", 
    x"698b", x"698a", x"6988", x"6986", x"6984", x"6982", x"6981", x"697f", 
    x"697d", x"697b", x"697a", x"6978", x"6976", x"6974", x"6972", x"6971", 
    x"696f", x"696d", x"696b", x"696a", x"6968", x"6966", x"6964", x"6962", 
    x"6961", x"695f", x"695d", x"695b", x"6959", x"6958", x"6956", x"6954", 
    x"6952", x"6951", x"694f", x"694d", x"694b", x"6949", x"6948", x"6946", 
    x"6944", x"6942", x"6940", x"693f", x"693d", x"693b", x"6939", x"6938", 
    x"6936", x"6934", x"6932", x"6930", x"692f", x"692d", x"692b", x"6929", 
    x"6927", x"6926", x"6924", x"6922", x"6920", x"691e", x"691d", x"691b", 
    x"6919", x"6917", x"6915", x"6914", x"6912", x"6910", x"690e", x"690d", 
    x"690b", x"6909", x"6907", x"6905", x"6904", x"6902", x"6900", x"68fe", 
    x"68fc", x"68fb", x"68f9", x"68f7", x"68f5", x"68f3", x"68f2", x"68f0", 
    x"68ee", x"68ec", x"68ea", x"68e9", x"68e7", x"68e5", x"68e3", x"68e1", 
    x"68e0", x"68de", x"68dc", x"68da", x"68d8", x"68d7", x"68d5", x"68d3", 
    x"68d1", x"68cf", x"68ce", x"68cc", x"68ca", x"68c8", x"68c6", x"68c5", 
    x"68c3", x"68c1", x"68bf", x"68bd", x"68bb", x"68ba", x"68b8", x"68b6", 
    x"68b4", x"68b2", x"68b1", x"68af", x"68ad", x"68ab", x"68a9", x"68a8", 
    x"68a6", x"68a4", x"68a2", x"68a0", x"689f", x"689d", x"689b", x"6899", 
    x"6897", x"6896", x"6894", x"6892", x"6890", x"688e", x"688c", x"688b", 
    x"6889", x"6887", x"6885", x"6883", x"6882", x"6880", x"687e", x"687c", 
    x"687a", x"6879", x"6877", x"6875", x"6873", x"6871", x"686f", x"686e", 
    x"686c", x"686a", x"6868", x"6866", x"6865", x"6863", x"6861", x"685f", 
    x"685d", x"685b", x"685a", x"6858", x"6856", x"6854", x"6852", x"6851", 
    x"684f", x"684d", x"684b", x"6849", x"6847", x"6846", x"6844", x"6842", 
    x"6840", x"683e", x"683c", x"683b", x"6839", x"6837", x"6835", x"6833", 
    x"6832", x"6830", x"682e", x"682c", x"682a", x"6828", x"6827", x"6825", 
    x"6823", x"6821", x"681f", x"681d", x"681c", x"681a", x"6818", x"6816", 
    x"6814", x"6812", x"6811", x"680f", x"680d", x"680b", x"6809", x"6807", 
    x"6806", x"6804", x"6802", x"6800", x"67fe", x"67fd", x"67fb", x"67f9", 
    x"67f7", x"67f5", x"67f3", x"67f2", x"67f0", x"67ee", x"67ec", x"67ea", 
    x"67e8", x"67e7", x"67e5", x"67e3", x"67e1", x"67df", x"67dd", x"67dc", 
    x"67da", x"67d8", x"67d6", x"67d4", x"67d2", x"67d0", x"67cf", x"67cd", 
    x"67cb", x"67c9", x"67c7", x"67c5", x"67c4", x"67c2", x"67c0", x"67be", 
    x"67bc", x"67ba", x"67b9", x"67b7", x"67b5", x"67b3", x"67b1", x"67af", 
    x"67ae", x"67ac", x"67aa", x"67a8", x"67a6", x"67a4", x"67a2", x"67a1", 
    x"679f", x"679d", x"679b", x"6799", x"6797", x"6796", x"6794", x"6792", 
    x"6790", x"678e", x"678c", x"678a", x"6789", x"6787", x"6785", x"6783", 
    x"6781", x"677f", x"677e", x"677c", x"677a", x"6778", x"6776", x"6774", 
    x"6772", x"6771", x"676f", x"676d", x"676b", x"6769", x"6767", x"6765", 
    x"6764", x"6762", x"6760", x"675e", x"675c", x"675a", x"6759", x"6757", 
    x"6755", x"6753", x"6751", x"674f", x"674d", x"674c", x"674a", x"6748", 
    x"6746", x"6744", x"6742", x"6740", x"673f", x"673d", x"673b", x"6739", 
    x"6737", x"6735", x"6733", x"6732", x"6730", x"672e", x"672c", x"672a", 
    x"6728", x"6726", x"6725", x"6723", x"6721", x"671f", x"671d", x"671b", 
    x"6719", x"6718", x"6716", x"6714", x"6712", x"6710", x"670e", x"670c", 
    x"670a", x"6709", x"6707", x"6705", x"6703", x"6701", x"66ff", x"66fd", 
    x"66fc", x"66fa", x"66f8", x"66f6", x"66f4", x"66f2", x"66f0", x"66ee", 
    x"66ed", x"66eb", x"66e9", x"66e7", x"66e5", x"66e3", x"66e1", x"66e0", 
    x"66de", x"66dc", x"66da", x"66d8", x"66d6", x"66d4", x"66d2", x"66d1", 
    x"66cf", x"66cd", x"66cb", x"66c9", x"66c7", x"66c5", x"66c3", x"66c2", 
    x"66c0", x"66be", x"66bc", x"66ba", x"66b8", x"66b6", x"66b4", x"66b3", 
    x"66b1", x"66af", x"66ad", x"66ab", x"66a9", x"66a7", x"66a5", x"66a4", 
    x"66a2", x"66a0", x"669e", x"669c", x"669a", x"6698", x"6696", x"6695", 
    x"6693", x"6691", x"668f", x"668d", x"668b", x"6689", x"6687", x"6686", 
    x"6684", x"6682", x"6680", x"667e", x"667c", x"667a", x"6678", x"6676", 
    x"6675", x"6673", x"6671", x"666f", x"666d", x"666b", x"6669", x"6667", 
    x"6666", x"6664", x"6662", x"6660", x"665e", x"665c", x"665a", x"6658", 
    x"6656", x"6655", x"6653", x"6651", x"664f", x"664d", x"664b", x"6649", 
    x"6647", x"6645", x"6644", x"6642", x"6640", x"663e", x"663c", x"663a", 
    x"6638", x"6636", x"6634", x"6633", x"6631", x"662f", x"662d", x"662b", 
    x"6629", x"6627", x"6625", x"6623", x"6622", x"6620", x"661e", x"661c", 
    x"661a", x"6618", x"6616", x"6614", x"6612", x"6610", x"660f", x"660d", 
    x"660b", x"6609", x"6607", x"6605", x"6603", x"6601", x"65ff", x"65fd", 
    x"65fc", x"65fa", x"65f8", x"65f6", x"65f4", x"65f2", x"65f0", x"65ee", 
    x"65ec", x"65ea", x"65e9", x"65e7", x"65e5", x"65e3", x"65e1", x"65df", 
    x"65dd", x"65db", x"65d9", x"65d7", x"65d6", x"65d4", x"65d2", x"65d0", 
    x"65ce", x"65cc", x"65ca", x"65c8", x"65c6", x"65c4", x"65c3", x"65c1", 
    x"65bf", x"65bd", x"65bb", x"65b9", x"65b7", x"65b5", x"65b3", x"65b1", 
    x"65af", x"65ae", x"65ac", x"65aa", x"65a8", x"65a6", x"65a4", x"65a2", 
    x"65a0", x"659e", x"659c", x"659a", x"6599", x"6597", x"6595", x"6593", 
    x"6591", x"658f", x"658d", x"658b", x"6589", x"6587", x"6585", x"6584", 
    x"6582", x"6580", x"657e", x"657c", x"657a", x"6578", x"6576", x"6574", 
    x"6572", x"6570", x"656e", x"656d", x"656b", x"6569", x"6567", x"6565", 
    x"6563", x"6561", x"655f", x"655d", x"655b", x"6559", x"6557", x"6556", 
    x"6554", x"6552", x"6550", x"654e", x"654c", x"654a", x"6548", x"6546", 
    x"6544", x"6542", x"6540", x"653e", x"653d", x"653b", x"6539", x"6537", 
    x"6535", x"6533", x"6531", x"652f", x"652d", x"652b", x"6529", x"6527", 
    x"6525", x"6524", x"6522", x"6520", x"651e", x"651c", x"651a", x"6518", 
    x"6516", x"6514", x"6512", x"6510", x"650e", x"650c", x"650a", x"6509", 
    x"6507", x"6505", x"6503", x"6501", x"64ff", x"64fd", x"64fb", x"64f9", 
    x"64f7", x"64f5", x"64f3", x"64f1", x"64ef", x"64ee", x"64ec", x"64ea", 
    x"64e8", x"64e6", x"64e4", x"64e2", x"64e0", x"64de", x"64dc", x"64da", 
    x"64d8", x"64d6", x"64d4", x"64d2", x"64d1", x"64cf", x"64cd", x"64cb", 
    x"64c9", x"64c7", x"64c5", x"64c3", x"64c1", x"64bf", x"64bd", x"64bb", 
    x"64b9", x"64b7", x"64b5", x"64b3", x"64b2", x"64b0", x"64ae", x"64ac", 
    x"64aa", x"64a8", x"64a6", x"64a4", x"64a2", x"64a0", x"649e", x"649c", 
    x"649a", x"6498", x"6496", x"6494", x"6492", x"6491", x"648f", x"648d", 
    x"648b", x"6489", x"6487", x"6485", x"6483", x"6481", x"647f", x"647d", 
    x"647b", x"6479", x"6477", x"6475", x"6473", x"6471", x"646f", x"646e", 
    x"646c", x"646a", x"6468", x"6466", x"6464", x"6462", x"6460", x"645e", 
    x"645c", x"645a", x"6458", x"6456", x"6454", x"6452", x"6450", x"644e", 
    x"644c", x"644a", x"6448", x"6447", x"6445", x"6443", x"6441", x"643f", 
    x"643d", x"643b", x"6439", x"6437", x"6435", x"6433", x"6431", x"642f", 
    x"642d", x"642b", x"6429", x"6427", x"6425", x"6423", x"6421", x"641f", 
    x"641d", x"641c", x"641a", x"6418", x"6416", x"6414", x"6412", x"6410", 
    x"640e", x"640c", x"640a", x"6408", x"6406", x"6404", x"6402", x"6400", 
    x"63fe", x"63fc", x"63fa", x"63f8", x"63f6", x"63f4", x"63f2", x"63f0", 
    x"63ee", x"63ec", x"63ea", x"63e9", x"63e7", x"63e5", x"63e3", x"63e1", 
    x"63df", x"63dd", x"63db", x"63d9", x"63d7", x"63d5", x"63d3", x"63d1", 
    x"63cf", x"63cd", x"63cb", x"63c9", x"63c7", x"63c5", x"63c3", x"63c1", 
    x"63bf", x"63bd", x"63bb", x"63b9", x"63b7", x"63b5", x"63b3", x"63b1", 
    x"63af", x"63ae", x"63ac", x"63aa", x"63a8", x"63a6", x"63a4", x"63a2", 
    x"63a0", x"639e", x"639c", x"639a", x"6398", x"6396", x"6394", x"6392", 
    x"6390", x"638e", x"638c", x"638a", x"6388", x"6386", x"6384", x"6382", 
    x"6380", x"637e", x"637c", x"637a", x"6378", x"6376", x"6374", x"6372", 
    x"6370", x"636e", x"636c", x"636a", x"6368", x"6366", x"6364", x"6362", 
    x"6360", x"635e", x"635d", x"635b", x"6359", x"6357", x"6355", x"6353", 
    x"6351", x"634f", x"634d", x"634b", x"6349", x"6347", x"6345", x"6343", 
    x"6341", x"633f", x"633d", x"633b", x"6339", x"6337", x"6335", x"6333", 
    x"6331", x"632f", x"632d", x"632b", x"6329", x"6327", x"6325", x"6323", 
    x"6321", x"631f", x"631d", x"631b", x"6319", x"6317", x"6315", x"6313", 
    x"6311", x"630f", x"630d", x"630b", x"6309", x"6307", x"6305", x"6303", 
    x"6301", x"62ff", x"62fd", x"62fb", x"62f9", x"62f7", x"62f5", x"62f3", 
    x"62f1", x"62ef", x"62ed", x"62eb", x"62e9", x"62e7", x"62e5", x"62e3", 
    x"62e1", x"62df", x"62dd", x"62db", x"62d9", x"62d7", x"62d5", x"62d3", 
    x"62d1", x"62cf", x"62cd", x"62cb", x"62c9", x"62c7", x"62c5", x"62c3", 
    x"62c1", x"62bf", x"62bd", x"62bb", x"62b9", x"62b7", x"62b5", x"62b3", 
    x"62b1", x"62af", x"62ad", x"62ab", x"62a9", x"62a7", x"62a5", x"62a3", 
    x"62a1", x"629f", x"629d", x"629b", x"6299", x"6297", x"6295", x"6293", 
    x"6291", x"628f", x"628d", x"628b", x"6289", x"6287", x"6285", x"6283", 
    x"6281", x"627f", x"627d", x"627b", x"6279", x"6277", x"6275", x"6273", 
    x"6271", x"626f", x"626d", x"626b", x"6269", x"6267", x"6265", x"6263", 
    x"6261", x"625f", x"625d", x"625b", x"6259", x"6257", x"6255", x"6253", 
    x"6251", x"624f", x"624d", x"624b", x"6249", x"6247", x"6245", x"6243", 
    x"6241", x"623f", x"623d", x"623b", x"6239", x"6237", x"6235", x"6233", 
    x"6231", x"622f", x"622d", x"622b", x"6229", x"6227", x"6225", x"6223", 
    x"6221", x"621f", x"621d", x"621b", x"6219", x"6217", x"6215", x"6213", 
    x"6211", x"620f", x"620d", x"620b", x"6208", x"6206", x"6204", x"6202", 
    x"6200", x"61fe", x"61fc", x"61fa", x"61f8", x"61f6", x"61f4", x"61f2", 
    x"61f0", x"61ee", x"61ec", x"61ea", x"61e8", x"61e6", x"61e4", x"61e2", 
    x"61e0", x"61de", x"61dc", x"61da", x"61d8", x"61d6", x"61d4", x"61d2", 
    x"61d0", x"61ce", x"61cc", x"61ca", x"61c8", x"61c6", x"61c4", x"61c2", 
    x"61c0", x"61be", x"61bc", x"61ba", x"61b8", x"61b5", x"61b3", x"61b1", 
    x"61af", x"61ad", x"61ab", x"61a9", x"61a7", x"61a5", x"61a3", x"61a1", 
    x"619f", x"619d", x"619b", x"6199", x"6197", x"6195", x"6193", x"6191", 
    x"618f", x"618d", x"618b", x"6189", x"6187", x"6185", x"6183", x"6181", 
    x"617f", x"617d", x"617b", x"6179", x"6176", x"6174", x"6172", x"6170", 
    x"616e", x"616c", x"616a", x"6168", x"6166", x"6164", x"6162", x"6160", 
    x"615e", x"615c", x"615a", x"6158", x"6156", x"6154", x"6152", x"6150", 
    x"614e", x"614c", x"614a", x"6148", x"6146", x"6143", x"6141", x"613f", 
    x"613d", x"613b", x"6139", x"6137", x"6135", x"6133", x"6131", x"612f", 
    x"612d", x"612b", x"6129", x"6127", x"6125", x"6123", x"6121", x"611f", 
    x"611d", x"611b", x"6119", x"6117", x"6114", x"6112", x"6110", x"610e", 
    x"610c", x"610a", x"6108", x"6106", x"6104", x"6102", x"6100", x"60fe", 
    x"60fc", x"60fa", x"60f8", x"60f6", x"60f4", x"60f2", x"60f0", x"60ee", 
    x"60eb", x"60e9", x"60e7", x"60e5", x"60e3", x"60e1", x"60df", x"60dd", 
    x"60db", x"60d9", x"60d7", x"60d5", x"60d3", x"60d1", x"60cf", x"60cd", 
    x"60cb", x"60c9", x"60c6", x"60c4", x"60c2", x"60c0", x"60be", x"60bc", 
    x"60ba", x"60b8", x"60b6", x"60b4", x"60b2", x"60b0", x"60ae", x"60ac", 
    x"60aa", x"60a8", x"60a6", x"60a4", x"60a1", x"609f", x"609d", x"609b", 
    x"6099", x"6097", x"6095", x"6093", x"6091", x"608f", x"608d", x"608b", 
    x"6089", x"6087", x"6085", x"6083", x"6080", x"607e", x"607c", x"607a", 
    x"6078", x"6076", x"6074", x"6072", x"6070", x"606e", x"606c", x"606a", 
    x"6068", x"6066", x"6064", x"6061", x"605f", x"605d", x"605b", x"6059", 
    x"6057", x"6055", x"6053", x"6051", x"604f", x"604d", x"604b", x"6049", 
    x"6047", x"6045", x"6042", x"6040", x"603e", x"603c", x"603a", x"6038", 
    x"6036", x"6034", x"6032", x"6030", x"602e", x"602c", x"602a", x"6028", 
    x"6025", x"6023", x"6021", x"601f", x"601d", x"601b", x"6019", x"6017", 
    x"6015", x"6013", x"6011", x"600f", x"600d", x"600a", x"6008", x"6006", 
    x"6004", x"6002", x"6000", x"5ffe", x"5ffc", x"5ffa", x"5ff8", x"5ff6", 
    x"5ff4", x"5ff2", x"5fef", x"5fed", x"5feb", x"5fe9", x"5fe7", x"5fe5", 
    x"5fe3", x"5fe1", x"5fdf", x"5fdd", x"5fdb", x"5fd9", x"5fd6", x"5fd4", 
    x"5fd2", x"5fd0", x"5fce", x"5fcc", x"5fca", x"5fc8", x"5fc6", x"5fc4", 
    x"5fc2", x"5fc0", x"5fbd", x"5fbb", x"5fb9", x"5fb7", x"5fb5", x"5fb3", 
    x"5fb1", x"5faf", x"5fad", x"5fab", x"5fa9", x"5fa7", x"5fa4", x"5fa2", 
    x"5fa0", x"5f9e", x"5f9c", x"5f9a", x"5f98", x"5f96", x"5f94", x"5f92", 
    x"5f90", x"5f8d", x"5f8b", x"5f89", x"5f87", x"5f85", x"5f83", x"5f81", 
    x"5f7f", x"5f7d", x"5f7b", x"5f79", x"5f76", x"5f74", x"5f72", x"5f70", 
    x"5f6e", x"5f6c", x"5f6a", x"5f68", x"5f66", x"5f64", x"5f61", x"5f5f", 
    x"5f5d", x"5f5b", x"5f59", x"5f57", x"5f55", x"5f53", x"5f51", x"5f4f", 
    x"5f4d", x"5f4a", x"5f48", x"5f46", x"5f44", x"5f42", x"5f40", x"5f3e", 
    x"5f3c", x"5f3a", x"5f38", x"5f35", x"5f33", x"5f31", x"5f2f", x"5f2d", 
    x"5f2b", x"5f29", x"5f27", x"5f25", x"5f23", x"5f20", x"5f1e", x"5f1c", 
    x"5f1a", x"5f18", x"5f16", x"5f14", x"5f12", x"5f10", x"5f0e", x"5f0b", 
    x"5f09", x"5f07", x"5f05", x"5f03", x"5f01", x"5eff", x"5efd", x"5efb", 
    x"5ef8", x"5ef6", x"5ef4", x"5ef2", x"5ef0", x"5eee", x"5eec", x"5eea", 
    x"5ee8", x"5ee6", x"5ee3", x"5ee1", x"5edf", x"5edd", x"5edb", x"5ed9", 
    x"5ed7", x"5ed5", x"5ed3", x"5ed0", x"5ece", x"5ecc", x"5eca", x"5ec8", 
    x"5ec6", x"5ec4", x"5ec2", x"5ec0", x"5ebd", x"5ebb", x"5eb9", x"5eb7", 
    x"5eb5", x"5eb3", x"5eb1", x"5eaf", x"5ead", x"5eaa", x"5ea8", x"5ea6", 
    x"5ea4", x"5ea2", x"5ea0", x"5e9e", x"5e9c", x"5e99", x"5e97", x"5e95", 
    x"5e93", x"5e91", x"5e8f", x"5e8d", x"5e8b", x"5e89", x"5e86", x"5e84", 
    x"5e82", x"5e80", x"5e7e", x"5e7c", x"5e7a", x"5e78", x"5e75", x"5e73", 
    x"5e71", x"5e6f", x"5e6d", x"5e6b", x"5e69", x"5e67", x"5e64", x"5e62", 
    x"5e60", x"5e5e", x"5e5c", x"5e5a", x"5e58", x"5e56", x"5e54", x"5e51", 
    x"5e4f", x"5e4d", x"5e4b", x"5e49", x"5e47", x"5e45", x"5e43", x"5e40", 
    x"5e3e", x"5e3c", x"5e3a", x"5e38", x"5e36", x"5e34", x"5e32", x"5e2f", 
    x"5e2d", x"5e2b", x"5e29", x"5e27", x"5e25", x"5e23", x"5e20", x"5e1e", 
    x"5e1c", x"5e1a", x"5e18", x"5e16", x"5e14", x"5e12", x"5e0f", x"5e0d", 
    x"5e0b", x"5e09", x"5e07", x"5e05", x"5e03", x"5e01", x"5dfe", x"5dfc", 
    x"5dfa", x"5df8", x"5df6", x"5df4", x"5df2", x"5def", x"5ded", x"5deb", 
    x"5de9", x"5de7", x"5de5", x"5de3", x"5de1", x"5dde", x"5ddc", x"5dda", 
    x"5dd8", x"5dd6", x"5dd4", x"5dd2", x"5dcf", x"5dcd", x"5dcb", x"5dc9", 
    x"5dc7", x"5dc5", x"5dc3", x"5dc0", x"5dbe", x"5dbc", x"5dba", x"5db8", 
    x"5db6", x"5db4", x"5db1", x"5daf", x"5dad", x"5dab", x"5da9", x"5da7", 
    x"5da5", x"5da3", x"5da0", x"5d9e", x"5d9c", x"5d9a", x"5d98", x"5d96", 
    x"5d94", x"5d91", x"5d8f", x"5d8d", x"5d8b", x"5d89", x"5d87", x"5d84", 
    x"5d82", x"5d80", x"5d7e", x"5d7c", x"5d7a", x"5d78", x"5d75", x"5d73", 
    x"5d71", x"5d6f", x"5d6d", x"5d6b", x"5d69", x"5d66", x"5d64", x"5d62", 
    x"5d60", x"5d5e", x"5d5c", x"5d5a", x"5d57", x"5d55", x"5d53", x"5d51", 
    x"5d4f", x"5d4d", x"5d4b", x"5d48", x"5d46", x"5d44", x"5d42", x"5d40", 
    x"5d3e", x"5d3b", x"5d39", x"5d37", x"5d35", x"5d33", x"5d31", x"5d2f", 
    x"5d2c", x"5d2a", x"5d28", x"5d26", x"5d24", x"5d22", x"5d1f", x"5d1d", 
    x"5d1b", x"5d19", x"5d17", x"5d15", x"5d13", x"5d10", x"5d0e", x"5d0c", 
    x"5d0a", x"5d08", x"5d06", x"5d03", x"5d01", x"5cff", x"5cfd", x"5cfb", 
    x"5cf9", x"5cf6", x"5cf4", x"5cf2", x"5cf0", x"5cee", x"5cec", x"5ce9", 
    x"5ce7", x"5ce5", x"5ce3", x"5ce1", x"5cdf", x"5cdd", x"5cda", x"5cd8", 
    x"5cd6", x"5cd4", x"5cd2", x"5cd0", x"5ccd", x"5ccb", x"5cc9", x"5cc7", 
    x"5cc5", x"5cc3", x"5cc0", x"5cbe", x"5cbc", x"5cba", x"5cb8", x"5cb6", 
    x"5cb3", x"5cb1", x"5caf", x"5cad", x"5cab", x"5ca9", x"5ca6", x"5ca4", 
    x"5ca2", x"5ca0", x"5c9e", x"5c9c", x"5c99", x"5c97", x"5c95", x"5c93", 
    x"5c91", x"5c8f", x"5c8c", x"5c8a", x"5c88", x"5c86", x"5c84", x"5c82", 
    x"5c7f", x"5c7d", x"5c7b", x"5c79", x"5c77", x"5c74", x"5c72", x"5c70", 
    x"5c6e", x"5c6c", x"5c6a", x"5c67", x"5c65", x"5c63", x"5c61", x"5c5f", 
    x"5c5d", x"5c5a", x"5c58", x"5c56", x"5c54", x"5c52", x"5c50", x"5c4d", 
    x"5c4b", x"5c49", x"5c47", x"5c45", x"5c42", x"5c40", x"5c3e", x"5c3c", 
    x"5c3a", x"5c38", x"5c35", x"5c33", x"5c31", x"5c2f", x"5c2d", x"5c2b", 
    x"5c28", x"5c26", x"5c24", x"5c22", x"5c20", x"5c1d", x"5c1b", x"5c19", 
    x"5c17", x"5c15", x"5c13", x"5c10", x"5c0e", x"5c0c", x"5c0a", x"5c08", 
    x"5c05", x"5c03", x"5c01", x"5bff", x"5bfd", x"5bfa", x"5bf8", x"5bf6", 
    x"5bf4", x"5bf2", x"5bf0", x"5bed", x"5beb", x"5be9", x"5be7", x"5be5", 
    x"5be2", x"5be0", x"5bde", x"5bdc", x"5bda", x"5bd8", x"5bd5", x"5bd3", 
    x"5bd1", x"5bcf", x"5bcd", x"5bca", x"5bc8", x"5bc6", x"5bc4", x"5bc2", 
    x"5bbf", x"5bbd", x"5bbb", x"5bb9", x"5bb7", x"5bb4", x"5bb2", x"5bb0", 
    x"5bae", x"5bac", x"5baa", x"5ba7", x"5ba5", x"5ba3", x"5ba1", x"5b9f", 
    x"5b9c", x"5b9a", x"5b98", x"5b96", x"5b94", x"5b91", x"5b8f", x"5b8d", 
    x"5b8b", x"5b89", x"5b86", x"5b84", x"5b82", x"5b80", x"5b7e", x"5b7b", 
    x"5b79", x"5b77", x"5b75", x"5b73", x"5b70", x"5b6e", x"5b6c", x"5b6a", 
    x"5b68", x"5b65", x"5b63", x"5b61", x"5b5f", x"5b5d", x"5b5a", x"5b58", 
    x"5b56", x"5b54", x"5b52", x"5b4f", x"5b4d", x"5b4b", x"5b49", x"5b47", 
    x"5b44", x"5b42", x"5b40", x"5b3e", x"5b3c", x"5b39", x"5b37", x"5b35", 
    x"5b33", x"5b31", x"5b2e", x"5b2c", x"5b2a", x"5b28", x"5b26", x"5b23", 
    x"5b21", x"5b1f", x"5b1d", x"5b1b", x"5b18", x"5b16", x"5b14", x"5b12", 
    x"5b0f", x"5b0d", x"5b0b", x"5b09", x"5b07", x"5b04", x"5b02", x"5b00", 
    x"5afe", x"5afc", x"5af9", x"5af7", x"5af5", x"5af3", x"5af1", x"5aee", 
    x"5aec", x"5aea", x"5ae8", x"5ae6", x"5ae3", x"5ae1", x"5adf", x"5add", 
    x"5ada", x"5ad8", x"5ad6", x"5ad4", x"5ad2", x"5acf", x"5acd", x"5acb", 
    x"5ac9", x"5ac7", x"5ac4", x"5ac2", x"5ac0", x"5abe", x"5abb", x"5ab9", 
    x"5ab7", x"5ab5", x"5ab3", x"5ab0", x"5aae", x"5aac", x"5aaa", x"5aa8", 
    x"5aa5", x"5aa3", x"5aa1", x"5a9f", x"5a9c", x"5a9a", x"5a98", x"5a96", 
    x"5a94", x"5a91", x"5a8f", x"5a8d", x"5a8b", x"5a88", x"5a86", x"5a84", 
    x"5a82", x"5a80", x"5a7d", x"5a7b", x"5a79", x"5a77", x"5a74", x"5a72", 
    x"5a70", x"5a6e", x"5a6c", x"5a69", x"5a67", x"5a65", x"5a63", x"5a60", 
    x"5a5e", x"5a5c", x"5a5a", x"5a58", x"5a55", x"5a53", x"5a51", x"5a4f", 
    x"5a4c", x"5a4a", x"5a48", x"5a46", x"5a43", x"5a41", x"5a3f", x"5a3d", 
    x"5a3b", x"5a38", x"5a36", x"5a34", x"5a32", x"5a2f", x"5a2d", x"5a2b", 
    x"5a29", x"5a27", x"5a24", x"5a22", x"5a20", x"5a1e", x"5a1b", x"5a19", 
    x"5a17", x"5a15", x"5a12", x"5a10", x"5a0e", x"5a0c", x"5a0a", x"5a07", 
    x"5a05", x"5a03", x"5a01", x"59fe", x"59fc", x"59fa", x"59f8", x"59f5", 
    x"59f3", x"59f1", x"59ef", x"59ec", x"59ea", x"59e8", x"59e6", x"59e4", 
    x"59e1", x"59df", x"59dd", x"59db", x"59d8", x"59d6", x"59d4", x"59d2", 
    x"59cf", x"59cd", x"59cb", x"59c9", x"59c6", x"59c4", x"59c2", x"59c0", 
    x"59bd", x"59bb", x"59b9", x"59b7", x"59b5", x"59b2", x"59b0", x"59ae", 
    x"59ac", x"59a9", x"59a7", x"59a5", x"59a3", x"59a0", x"599e", x"599c", 
    x"599a", x"5997", x"5995", x"5993", x"5991", x"598e", x"598c", x"598a", 
    x"5988", x"5985", x"5983", x"5981", x"597f", x"597c", x"597a", x"5978", 
    x"5976", x"5973", x"5971", x"596f", x"596d", x"596a", x"5968", x"5966", 
    x"5964", x"5961", x"595f", x"595d", x"595b", x"5958", x"5956", x"5954", 
    x"5952", x"594f", x"594d", x"594b", x"5949", x"5946", x"5944", x"5942", 
    x"5940", x"593d", x"593b", x"5939", x"5937", x"5934", x"5932", x"5930", 
    x"592e", x"592b", x"5929", x"5927", x"5925", x"5922", x"5920", x"591e", 
    x"591c", x"5919", x"5917", x"5915", x"5913", x"5910", x"590e", x"590c", 
    x"590a", x"5907", x"5905", x"5903", x"5901", x"58fe", x"58fc", x"58fa", 
    x"58f8", x"58f5", x"58f3", x"58f1", x"58ee", x"58ec", x"58ea", x"58e8", 
    x"58e5", x"58e3", x"58e1", x"58df", x"58dc", x"58da", x"58d8", x"58d6", 
    x"58d3", x"58d1", x"58cf", x"58cd", x"58ca", x"58c8", x"58c6", x"58c4", 
    x"58c1", x"58bf", x"58bd", x"58ba", x"58b8", x"58b6", x"58b4", x"58b1", 
    x"58af", x"58ad", x"58ab", x"58a8", x"58a6", x"58a4", x"58a2", x"589f", 
    x"589d", x"589b", x"5898", x"5896", x"5894", x"5892", x"588f", x"588d", 
    x"588b", x"5889", x"5886", x"5884", x"5882", x"5880", x"587d", x"587b", 
    x"5879", x"5876", x"5874", x"5872", x"5870", x"586d", x"586b", x"5869", 
    x"5867", x"5864", x"5862", x"5860", x"585d", x"585b", x"5859", x"5857", 
    x"5854", x"5852", x"5850", x"584e", x"584b", x"5849", x"5847", x"5844", 
    x"5842", x"5840", x"583e", x"583b", x"5839", x"5837", x"5835", x"5832", 
    x"5830", x"582e", x"582b", x"5829", x"5827", x"5825", x"5822", x"5820", 
    x"581e", x"581b", x"5819", x"5817", x"5815", x"5812", x"5810", x"580e", 
    x"580c", x"5809", x"5807", x"5805", x"5802", x"5800", x"57fe", x"57fc", 
    x"57f9", x"57f7", x"57f5", x"57f2", x"57f0", x"57ee", x"57ec", x"57e9", 
    x"57e7", x"57e5", x"57e2", x"57e0", x"57de", x"57dc", x"57d9", x"57d7", 
    x"57d5", x"57d2", x"57d0", x"57ce", x"57cc", x"57c9", x"57c7", x"57c5", 
    x"57c2", x"57c0", x"57be", x"57bc", x"57b9", x"57b7", x"57b5", x"57b2", 
    x"57b0", x"57ae", x"57ac", x"57a9", x"57a7", x"57a5", x"57a2", x"57a0", 
    x"579e", x"579c", x"5799", x"5797", x"5795", x"5792", x"5790", x"578e", 
    x"578b", x"5789", x"5787", x"5785", x"5782", x"5780", x"577e", x"577b", 
    x"5779", x"5777", x"5775", x"5772", x"5770", x"576e", x"576b", x"5769", 
    x"5767", x"5765", x"5762", x"5760", x"575e", x"575b", x"5759", x"5757", 
    x"5754", x"5752", x"5750", x"574e", x"574b", x"5749", x"5747", x"5744", 
    x"5742", x"5740", x"573d", x"573b", x"5739", x"5737", x"5734", x"5732", 
    x"5730", x"572d", x"572b", x"5729", x"5726", x"5724", x"5722", x"5720", 
    x"571d", x"571b", x"5719", x"5716", x"5714", x"5712", x"570f", x"570d", 
    x"570b", x"5709", x"5706", x"5704", x"5702", x"56ff", x"56fd", x"56fb", 
    x"56f8", x"56f6", x"56f4", x"56f1", x"56ef", x"56ed", x"56eb", x"56e8", 
    x"56e6", x"56e4", x"56e1", x"56df", x"56dd", x"56da", x"56d8", x"56d6", 
    x"56d3", x"56d1", x"56cf", x"56cd", x"56ca", x"56c8", x"56c6", x"56c3", 
    x"56c1", x"56bf", x"56bc", x"56ba", x"56b8", x"56b5", x"56b3", x"56b1", 
    x"56af", x"56ac", x"56aa", x"56a8", x"56a5", x"56a3", x"56a1", x"569e", 
    x"569c", x"569a", x"5697", x"5695", x"5693", x"5690", x"568e", x"568c", 
    x"568a", x"5687", x"5685", x"5683", x"5680", x"567e", x"567c", x"5679", 
    x"5677", x"5675", x"5672", x"5670", x"566e", x"566b", x"5669", x"5667", 
    x"5664", x"5662", x"5660", x"565e", x"565b", x"5659", x"5657", x"5654", 
    x"5652", x"5650", x"564d", x"564b", x"5649", x"5646", x"5644", x"5642", 
    x"563f", x"563d", x"563b", x"5638", x"5636", x"5634", x"5631", x"562f", 
    x"562d", x"562a", x"5628", x"5626", x"5623", x"5621", x"561f", x"561d", 
    x"561a", x"5618", x"5616", x"5613", x"5611", x"560f", x"560c", x"560a", 
    x"5608", x"5605", x"5603", x"5601", x"55fe", x"55fc", x"55fa", x"55f7", 
    x"55f5", x"55f3", x"55f0", x"55ee", x"55ec", x"55e9", x"55e7", x"55e5", 
    x"55e2", x"55e0", x"55de", x"55db", x"55d9", x"55d7", x"55d4", x"55d2", 
    x"55d0", x"55cd", x"55cb", x"55c9", x"55c6", x"55c4", x"55c2", x"55bf", 
    x"55bd", x"55bb", x"55b8", x"55b6", x"55b4", x"55b1", x"55af", x"55ad", 
    x"55aa", x"55a8", x"55a6", x"55a3", x"55a1", x"559f", x"559c", x"559a", 
    x"5598", x"5595", x"5593", x"5591", x"558e", x"558c", x"558a", x"5587", 
    x"5585", x"5583", x"5580", x"557e", x"557c", x"5579", x"5577", x"5575", 
    x"5572", x"5570", x"556e", x"556b", x"5569", x"5567", x"5564", x"5562", 
    x"5560", x"555d", x"555b", x"5559", x"5556", x"5554", x"5552", x"554f", 
    x"554d", x"554b", x"5548", x"5546", x"5543", x"5541", x"553f", x"553c", 
    x"553a", x"5538", x"5535", x"5533", x"5531", x"552e", x"552c", x"552a", 
    x"5527", x"5525", x"5523", x"5520", x"551e", x"551c", x"5519", x"5517", 
    x"5515", x"5512", x"5510", x"550e", x"550b", x"5509", x"5506", x"5504", 
    x"5502", x"54ff", x"54fd", x"54fb", x"54f8", x"54f6", x"54f4", x"54f1", 
    x"54ef", x"54ed", x"54ea", x"54e8", x"54e6", x"54e3", x"54e1", x"54df", 
    x"54dc", x"54da", x"54d7", x"54d5", x"54d3", x"54d0", x"54ce", x"54cc", 
    x"54c9", x"54c7", x"54c5", x"54c2", x"54c0", x"54be", x"54bb", x"54b9", 
    x"54b7", x"54b4", x"54b2", x"54af", x"54ad", x"54ab", x"54a8", x"54a6", 
    x"54a4", x"54a1", x"549f", x"549d", x"549a", x"5498", x"5496", x"5493", 
    x"5491", x"548e", x"548c", x"548a", x"5487", x"5485", x"5483", x"5480", 
    x"547e", x"547c", x"5479", x"5477", x"5475", x"5472", x"5470", x"546d", 
    x"546b", x"5469", x"5466", x"5464", x"5462", x"545f", x"545d", x"545b", 
    x"5458", x"5456", x"5453", x"5451", x"544f", x"544c", x"544a", x"5448", 
    x"5445", x"5443", x"5441", x"543e", x"543c", x"5439", x"5437", x"5435", 
    x"5432", x"5430", x"542e", x"542b", x"5429", x"5427", x"5424", x"5422", 
    x"541f", x"541d", x"541b", x"5418", x"5416", x"5414", x"5411", x"540f", 
    x"540c", x"540a", x"5408", x"5405", x"5403", x"5401", x"53fe", x"53fc", 
    x"53fa", x"53f7", x"53f5", x"53f2", x"53f0", x"53ee", x"53eb", x"53e9", 
    x"53e7", x"53e4", x"53e2", x"53df", x"53dd", x"53db", x"53d8", x"53d6", 
    x"53d4", x"53d1", x"53cf", x"53cc", x"53ca", x"53c8", x"53c5", x"53c3", 
    x"53c1", x"53be", x"53bc", x"53b9", x"53b7", x"53b5", x"53b2", x"53b0", 
    x"53ae", x"53ab", x"53a9", x"53a6", x"53a4", x"53a2", x"539f", x"539d", 
    x"539b", x"5398", x"5396", x"5393", x"5391", x"538f", x"538c", x"538a", 
    x"5387", x"5385", x"5383", x"5380", x"537e", x"537c", x"5379", x"5377", 
    x"5374", x"5372", x"5370", x"536d", x"536b", x"5369", x"5366", x"5364", 
    x"5361", x"535f", x"535d", x"535a", x"5358", x"5355", x"5353", x"5351", 
    x"534e", x"534c", x"534a", x"5347", x"5345", x"5342", x"5340", x"533e", 
    x"533b", x"5339", x"5336", x"5334", x"5332", x"532f", x"532d", x"532a", 
    x"5328", x"5326", x"5323", x"5321", x"531f", x"531c", x"531a", x"5317", 
    x"5315", x"5313", x"5310", x"530e", x"530b", x"5309", x"5307", x"5304", 
    x"5302", x"52ff", x"52fd", x"52fb", x"52f8", x"52f6", x"52f4", x"52f1", 
    x"52ef", x"52ec", x"52ea", x"52e8", x"52e5", x"52e3", x"52e0", x"52de", 
    x"52dc", x"52d9", x"52d7", x"52d4", x"52d2", x"52d0", x"52cd", x"52cb", 
    x"52c8", x"52c6", x"52c4", x"52c1", x"52bf", x"52bc", x"52ba", x"52b8", 
    x"52b5", x"52b3", x"52b0", x"52ae", x"52ac", x"52a9", x"52a7", x"52a4", 
    x"52a2", x"52a0", x"529d", x"529b", x"5298", x"5296", x"5294", x"5291", 
    x"528f", x"528c", x"528a", x"5288", x"5285", x"5283", x"5280", x"527e", 
    x"527c", x"5279", x"5277", x"5274", x"5272", x"5270", x"526d", x"526b", 
    x"5268", x"5266", x"5264", x"5261", x"525f", x"525c", x"525a", x"5258", 
    x"5255", x"5253", x"5250", x"524e", x"524c", x"5249", x"5247", x"5244", 
    x"5242", x"5240", x"523d", x"523b", x"5238", x"5236", x"5233", x"5231", 
    x"522f", x"522c", x"522a", x"5227", x"5225", x"5223", x"5220", x"521e", 
    x"521b", x"5219", x"5217", x"5214", x"5212", x"520f", x"520d", x"520b", 
    x"5208", x"5206", x"5203", x"5201", x"51fe", x"51fc", x"51fa", x"51f7", 
    x"51f5", x"51f2", x"51f0", x"51ee", x"51eb", x"51e9", x"51e6", x"51e4", 
    x"51e2", x"51df", x"51dd", x"51da", x"51d8", x"51d5", x"51d3", x"51d1", 
    x"51ce", x"51cc", x"51c9", x"51c7", x"51c5", x"51c2", x"51c0", x"51bd", 
    x"51bb", x"51b8", x"51b6", x"51b4", x"51b1", x"51af", x"51ac", x"51aa", 
    x"51a8", x"51a5", x"51a3", x"51a0", x"519e", x"519b", x"5199", x"5197", 
    x"5194", x"5192", x"518f", x"518d", x"518a", x"5188", x"5186", x"5183", 
    x"5181", x"517e", x"517c", x"517a", x"5177", x"5175", x"5172", x"5170", 
    x"516d", x"516b", x"5169", x"5166", x"5164", x"5161", x"515f", x"515c", 
    x"515a", x"5158", x"5155", x"5153", x"5150", x"514e", x"514b", x"5149", 
    x"5147", x"5144", x"5142", x"513f", x"513d", x"513a", x"5138", x"5136", 
    x"5133", x"5131", x"512e", x"512c", x"5129", x"5127", x"5125", x"5122", 
    x"5120", x"511d", x"511b", x"5118", x"5116", x"5114", x"5111", x"510f", 
    x"510c", x"510a", x"5107", x"5105", x"5103", x"5100", x"50fe", x"50fb", 
    x"50f9", x"50f6", x"50f4", x"50f2", x"50ef", x"50ed", x"50ea", x"50e8", 
    x"50e5", x"50e3", x"50e0", x"50de", x"50dc", x"50d9", x"50d7", x"50d4", 
    x"50d2", x"50cf", x"50cd", x"50cb", x"50c8", x"50c6", x"50c3", x"50c1", 
    x"50be", x"50bc", x"50ba", x"50b7", x"50b5", x"50b2", x"50b0", x"50ad", 
    x"50ab", x"50a8", x"50a6", x"50a4", x"50a1", x"509f", x"509c", x"509a", 
    x"5097", x"5095", x"5092", x"5090", x"508e", x"508b", x"5089", x"5086", 
    x"5084", x"5081", x"507f", x"507c", x"507a", x"5078", x"5075", x"5073", 
    x"5070", x"506e", x"506b", x"5069", x"5067", x"5064", x"5062", x"505f", 
    x"505d", x"505a", x"5058", x"5055", x"5053", x"5050", x"504e", x"504c", 
    x"5049", x"5047", x"5044", x"5042", x"503f", x"503d", x"503a", x"5038", 
    x"5036", x"5033", x"5031", x"502e", x"502c", x"5029", x"5027", x"5024", 
    x"5022", x"5020", x"501d", x"501b", x"5018", x"5016", x"5013", x"5011", 
    x"500e", x"500c", x"5009", x"5007", x"5005", x"5002", x"5000", x"4ffd", 
    x"4ffb", x"4ff8", x"4ff6", x"4ff3", x"4ff1", x"4fef", x"4fec", x"4fea", 
    x"4fe7", x"4fe5", x"4fe2", x"4fe0", x"4fdd", x"4fdb", x"4fd8", x"4fd6", 
    x"4fd4", x"4fd1", x"4fcf", x"4fcc", x"4fca", x"4fc7", x"4fc5", x"4fc2", 
    x"4fc0", x"4fbd", x"4fbb", x"4fb8", x"4fb6", x"4fb4", x"4fb1", x"4faf", 
    x"4fac", x"4faa", x"4fa7", x"4fa5", x"4fa2", x"4fa0", x"4f9d", x"4f9b", 
    x"4f99", x"4f96", x"4f94", x"4f91", x"4f8f", x"4f8c", x"4f8a", x"4f87", 
    x"4f85", x"4f82", x"4f80", x"4f7d", x"4f7b", x"4f79", x"4f76", x"4f74", 
    x"4f71", x"4f6f", x"4f6c", x"4f6a", x"4f67", x"4f65", x"4f62", x"4f60", 
    x"4f5d", x"4f5b", x"4f58", x"4f56", x"4f54", x"4f51", x"4f4f", x"4f4c", 
    x"4f4a", x"4f47", x"4f45", x"4f42", x"4f40", x"4f3d", x"4f3b", x"4f38", 
    x"4f36", x"4f33", x"4f31", x"4f2f", x"4f2c", x"4f2a", x"4f27", x"4f25", 
    x"4f22", x"4f20", x"4f1d", x"4f1b", x"4f18", x"4f16", x"4f13", x"4f11", 
    x"4f0e", x"4f0c", x"4f0a", x"4f07", x"4f05", x"4f02", x"4f00", x"4efd", 
    x"4efb", x"4ef8", x"4ef6", x"4ef3", x"4ef1", x"4eee", x"4eec", x"4ee9", 
    x"4ee7", x"4ee4", x"4ee2", x"4edf", x"4edd", x"4edb", x"4ed8", x"4ed6", 
    x"4ed3", x"4ed1", x"4ece", x"4ecc", x"4ec9", x"4ec7", x"4ec4", x"4ec2", 
    x"4ebf", x"4ebd", x"4eba", x"4eb8", x"4eb5", x"4eb3", x"4eb0", x"4eae", 
    x"4eab", x"4ea9", x"4ea7", x"4ea4", x"4ea2", x"4e9f", x"4e9d", x"4e9a", 
    x"4e98", x"4e95", x"4e93", x"4e90", x"4e8e", x"4e8b", x"4e89", x"4e86", 
    x"4e84", x"4e81", x"4e7f", x"4e7c", x"4e7a", x"4e77", x"4e75", x"4e72", 
    x"4e70", x"4e6d", x"4e6b", x"4e68", x"4e66", x"4e64", x"4e61", x"4e5f", 
    x"4e5c", x"4e5a", x"4e57", x"4e55", x"4e52", x"4e50", x"4e4d", x"4e4b", 
    x"4e48", x"4e46", x"4e43", x"4e41", x"4e3e", x"4e3c", x"4e39", x"4e37", 
    x"4e34", x"4e32", x"4e2f", x"4e2d", x"4e2a", x"4e28", x"4e25", x"4e23", 
    x"4e20", x"4e1e", x"4e1b", x"4e19", x"4e16", x"4e14", x"4e11", x"4e0f", 
    x"4e0d", x"4e0a", x"4e08", x"4e05", x"4e03", x"4e00", x"4dfe", x"4dfb", 
    x"4df9", x"4df6", x"4df4", x"4df1", x"4def", x"4dec", x"4dea", x"4de7", 
    x"4de5", x"4de2", x"4de0", x"4ddd", x"4ddb", x"4dd8", x"4dd6", x"4dd3", 
    x"4dd1", x"4dce", x"4dcc", x"4dc9", x"4dc7", x"4dc4", x"4dc2", x"4dbf", 
    x"4dbd", x"4dba", x"4db8", x"4db5", x"4db3", x"4db0", x"4dae", x"4dab", 
    x"4da9", x"4da6", x"4da4", x"4da1", x"4d9f", x"4d9c", x"4d9a", x"4d97", 
    x"4d95", x"4d92", x"4d90", x"4d8d", x"4d8b", x"4d88", x"4d86", x"4d83", 
    x"4d81", x"4d7e", x"4d7c", x"4d79", x"4d77", x"4d74", x"4d72", x"4d6f", 
    x"4d6d", x"4d6a", x"4d68", x"4d65", x"4d63", x"4d60", x"4d5e", x"4d5b", 
    x"4d59", x"4d56", x"4d54", x"4d51", x"4d4f", x"4d4c", x"4d4a", x"4d47", 
    x"4d45", x"4d42", x"4d40", x"4d3d", x"4d3b", x"4d38", x"4d36", x"4d33", 
    x"4d31", x"4d2e", x"4d2c", x"4d29", x"4d27", x"4d24", x"4d22", x"4d1f", 
    x"4d1d", x"4d1a", x"4d18", x"4d15", x"4d13", x"4d10", x"4d0e", x"4d0b", 
    x"4d09", x"4d06", x"4d04", x"4d01", x"4cff", x"4cfc", x"4cfa", x"4cf7", 
    x"4cf4", x"4cf2", x"4cef", x"4ced", x"4cea", x"4ce8", x"4ce5", x"4ce3", 
    x"4ce0", x"4cde", x"4cdb", x"4cd9", x"4cd6", x"4cd4", x"4cd1", x"4ccf", 
    x"4ccc", x"4cca", x"4cc7", x"4cc5", x"4cc2", x"4cc0", x"4cbd", x"4cbb", 
    x"4cb8", x"4cb6", x"4cb3", x"4cb1", x"4cae", x"4cac", x"4ca9", x"4ca7", 
    x"4ca4", x"4ca2", x"4c9f", x"4c9d", x"4c9a", x"4c97", x"4c95", x"4c92", 
    x"4c90", x"4c8d", x"4c8b", x"4c88", x"4c86", x"4c83", x"4c81", x"4c7e", 
    x"4c7c", x"4c79", x"4c77", x"4c74", x"4c72", x"4c6f", x"4c6d", x"4c6a", 
    x"4c68", x"4c65", x"4c63", x"4c60", x"4c5e", x"4c5b", x"4c59", x"4c56", 
    x"4c53", x"4c51", x"4c4e", x"4c4c", x"4c49", x"4c47", x"4c44", x"4c42", 
    x"4c3f", x"4c3d", x"4c3a", x"4c38", x"4c35", x"4c33", x"4c30", x"4c2e", 
    x"4c2b", x"4c29", x"4c26", x"4c24", x"4c21", x"4c1e", x"4c1c", x"4c19", 
    x"4c17", x"4c14", x"4c12", x"4c0f", x"4c0d", x"4c0a", x"4c08", x"4c05", 
    x"4c03", x"4c00", x"4bfe", x"4bfb", x"4bf9", x"4bf6", x"4bf4", x"4bf1", 
    x"4bee", x"4bec", x"4be9", x"4be7", x"4be4", x"4be2", x"4bdf", x"4bdd", 
    x"4bda", x"4bd8", x"4bd5", x"4bd3", x"4bd0", x"4bce", x"4bcb", x"4bc8", 
    x"4bc6", x"4bc3", x"4bc1", x"4bbe", x"4bbc", x"4bb9", x"4bb7", x"4bb4", 
    x"4bb2", x"4baf", x"4bad", x"4baa", x"4ba8", x"4ba5", x"4ba2", x"4ba0", 
    x"4b9d", x"4b9b", x"4b98", x"4b96", x"4b93", x"4b91", x"4b8e", x"4b8c", 
    x"4b89", x"4b87", x"4b84", x"4b82", x"4b7f", x"4b7c", x"4b7a", x"4b77", 
    x"4b75", x"4b72", x"4b70", x"4b6d", x"4b6b", x"4b68", x"4b66", x"4b63", 
    x"4b61", x"4b5e", x"4b5b", x"4b59", x"4b56", x"4b54", x"4b51", x"4b4f", 
    x"4b4c", x"4b4a", x"4b47", x"4b45", x"4b42", x"4b40", x"4b3d", x"4b3a", 
    x"4b38", x"4b35", x"4b33", x"4b30", x"4b2e", x"4b2b", x"4b29", x"4b26", 
    x"4b24", x"4b21", x"4b1e", x"4b1c", x"4b19", x"4b17", x"4b14", x"4b12", 
    x"4b0f", x"4b0d", x"4b0a", x"4b08", x"4b05", x"4b02", x"4b00", x"4afd", 
    x"4afb", x"4af8", x"4af6", x"4af3", x"4af1", x"4aee", x"4aec", x"4ae9", 
    x"4ae6", x"4ae4", x"4ae1", x"4adf", x"4adc", x"4ada", x"4ad7", x"4ad5", 
    x"4ad2", x"4ad0", x"4acd", x"4aca", x"4ac8", x"4ac5", x"4ac3", x"4ac0", 
    x"4abe", x"4abb", x"4ab9", x"4ab6", x"4ab3", x"4ab1", x"4aae", x"4aac", 
    x"4aa9", x"4aa7", x"4aa4", x"4aa2", x"4a9f", x"4a9d", x"4a9a", x"4a97", 
    x"4a95", x"4a92", x"4a90", x"4a8d", x"4a8b", x"4a88", x"4a86", x"4a83", 
    x"4a80", x"4a7e", x"4a7b", x"4a79", x"4a76", x"4a74", x"4a71", x"4a6f", 
    x"4a6c", x"4a69", x"4a67", x"4a64", x"4a62", x"4a5f", x"4a5d", x"4a5a", 
    x"4a58", x"4a55", x"4a52", x"4a50", x"4a4d", x"4a4b", x"4a48", x"4a46", 
    x"4a43", x"4a41", x"4a3e", x"4a3b", x"4a39", x"4a36", x"4a34", x"4a31", 
    x"4a2f", x"4a2c", x"4a29", x"4a27", x"4a24", x"4a22", x"4a1f", x"4a1d", 
    x"4a1a", x"4a18", x"4a15", x"4a12", x"4a10", x"4a0d", x"4a0b", x"4a08", 
    x"4a06", x"4a03", x"4a00", x"49fe", x"49fb", x"49f9", x"49f6", x"49f4", 
    x"49f1", x"49ef", x"49ec", x"49e9", x"49e7", x"49e4", x"49e2", x"49df", 
    x"49dd", x"49da", x"49d7", x"49d5", x"49d2", x"49d0", x"49cd", x"49cb", 
    x"49c8", x"49c5", x"49c3", x"49c0", x"49be", x"49bb", x"49b9", x"49b6", 
    x"49b4", x"49b1", x"49ae", x"49ac", x"49a9", x"49a7", x"49a4", x"49a2", 
    x"499f", x"499c", x"499a", x"4997", x"4995", x"4992", x"4990", x"498d", 
    x"498a", x"4988", x"4985", x"4983", x"4980", x"497e", x"497b", x"4978", 
    x"4976", x"4973", x"4971", x"496e", x"496c", x"4969", x"4966", x"4964", 
    x"4961", x"495f", x"495c", x"495a", x"4957", x"4954", x"4952", x"494f", 
    x"494d", x"494a", x"4947", x"4945", x"4942", x"4940", x"493d", x"493b", 
    x"4938", x"4935", x"4933", x"4930", x"492e", x"492b", x"4929", x"4926", 
    x"4923", x"4921", x"491e", x"491c", x"4919", x"4917", x"4914", x"4911", 
    x"490f", x"490c", x"490a", x"4907", x"4904", x"4902", x"48ff", x"48fd", 
    x"48fa", x"48f8", x"48f5", x"48f2", x"48f0", x"48ed", x"48eb", x"48e8", 
    x"48e5", x"48e3", x"48e0", x"48de", x"48db", x"48d9", x"48d6", x"48d3", 
    x"48d1", x"48ce", x"48cc", x"48c9", x"48c6", x"48c4", x"48c1", x"48bf", 
    x"48bc", x"48ba", x"48b7", x"48b4", x"48b2", x"48af", x"48ad", x"48aa", 
    x"48a7", x"48a5", x"48a2", x"48a0", x"489d", x"489b", x"4898", x"4895", 
    x"4893", x"4890", x"488e", x"488b", x"4888", x"4886", x"4883", x"4881", 
    x"487e", x"487b", x"4879", x"4876", x"4874", x"4871", x"486f", x"486c", 
    x"4869", x"4867", x"4864", x"4862", x"485f", x"485c", x"485a", x"4857", 
    x"4855", x"4852", x"484f", x"484d", x"484a", x"4848", x"4845", x"4842", 
    x"4840", x"483d", x"483b", x"4838", x"4835", x"4833", x"4830", x"482e", 
    x"482b", x"4829", x"4826", x"4823", x"4821", x"481e", x"481c", x"4819", 
    x"4816", x"4814", x"4811", x"480f", x"480c", x"4809", x"4807", x"4804", 
    x"4802", x"47ff", x"47fc", x"47fa", x"47f7", x"47f5", x"47f2", x"47ef", 
    x"47ed", x"47ea", x"47e8", x"47e5", x"47e2", x"47e0", x"47dd", x"47db", 
    x"47d8", x"47d5", x"47d3", x"47d0", x"47ce", x"47cb", x"47c8", x"47c6", 
    x"47c3", x"47c1", x"47be", x"47bb", x"47b9", x"47b6", x"47b4", x"47b1", 
    x"47ae", x"47ac", x"47a9", x"47a7", x"47a4", x"47a1", x"479f", x"479c", 
    x"479a", x"4797", x"4794", x"4792", x"478f", x"478d", x"478a", x"4787", 
    x"4785", x"4782", x"4780", x"477d", x"477a", x"4778", x"4775", x"4772", 
    x"4770", x"476d", x"476b", x"4768", x"4765", x"4763", x"4760", x"475e", 
    x"475b", x"4758", x"4756", x"4753", x"4751", x"474e", x"474b", x"4749", 
    x"4746", x"4744", x"4741", x"473e", x"473c", x"4739", x"4736", x"4734", 
    x"4731", x"472f", x"472c", x"4729", x"4727", x"4724", x"4722", x"471f", 
    x"471c", x"471a", x"4717", x"4715", x"4712", x"470f", x"470d", x"470a", 
    x"4707", x"4705", x"4702", x"4700", x"46fd", x"46fa", x"46f8", x"46f5", 
    x"46f3", x"46f0", x"46ed", x"46eb", x"46e8", x"46e5", x"46e3", x"46e0", 
    x"46de", x"46db", x"46d8", x"46d6", x"46d3", x"46d1", x"46ce", x"46cb", 
    x"46c9", x"46c6", x"46c3", x"46c1", x"46be", x"46bc", x"46b9", x"46b6", 
    x"46b4", x"46b1", x"46af", x"46ac", x"46a9", x"46a7", x"46a4", x"46a1", 
    x"469f", x"469c", x"469a", x"4697", x"4694", x"4692", x"468f", x"468c", 
    x"468a", x"4687", x"4685", x"4682", x"467f", x"467d", x"467a", x"4677", 
    x"4675", x"4672", x"4670", x"466d", x"466a", x"4668", x"4665", x"4662", 
    x"4660", x"465d", x"465b", x"4658", x"4655", x"4653", x"4650", x"464d", 
    x"464b", x"4648", x"4646", x"4643", x"4640", x"463e", x"463b", x"4638", 
    x"4636", x"4633", x"4631", x"462e", x"462b", x"4629", x"4626", x"4623", 
    x"4621", x"461e", x"461c", x"4619", x"4616", x"4614", x"4611", x"460e", 
    x"460c", x"4609", x"4607", x"4604", x"4601", x"45ff", x"45fc", x"45f9", 
    x"45f7", x"45f4", x"45f2", x"45ef", x"45ec", x"45ea", x"45e7", x"45e4", 
    x"45e2", x"45df", x"45dc", x"45da", x"45d7", x"45d5", x"45d2", x"45cf", 
    x"45cd", x"45ca", x"45c7", x"45c5", x"45c2", x"45bf", x"45bd", x"45ba", 
    x"45b8", x"45b5", x"45b2", x"45b0", x"45ad", x"45aa", x"45a8", x"45a5", 
    x"45a3", x"45a0", x"459d", x"459b", x"4598", x"4595", x"4593", x"4590", 
    x"458d", x"458b", x"4588", x"4586", x"4583", x"4580", x"457e", x"457b", 
    x"4578", x"4576", x"4573", x"4570", x"456e", x"456b", x"4568", x"4566", 
    x"4563", x"4561", x"455e", x"455b", x"4559", x"4556", x"4553", x"4551", 
    x"454e", x"454b", x"4549", x"4546", x"4544", x"4541", x"453e", x"453c", 
    x"4539", x"4536", x"4534", x"4531", x"452e", x"452c", x"4529", x"4526", 
    x"4524", x"4521", x"451f", x"451c", x"4519", x"4517", x"4514", x"4511", 
    x"450f", x"450c", x"4509", x"4507", x"4504", x"4501", x"44ff", x"44fc", 
    x"44f9", x"44f7", x"44f4", x"44f2", x"44ef", x"44ec", x"44ea", x"44e7", 
    x"44e4", x"44e2", x"44df", x"44dc", x"44da", x"44d7", x"44d4", x"44d2", 
    x"44cf", x"44cc", x"44ca", x"44c7", x"44c5", x"44c2", x"44bf", x"44bd", 
    x"44ba", x"44b7", x"44b5", x"44b2", x"44af", x"44ad", x"44aa", x"44a7", 
    x"44a5", x"44a2", x"449f", x"449d", x"449a", x"4497", x"4495", x"4492", 
    x"448f", x"448d", x"448a", x"4488", x"4485", x"4482", x"4480", x"447d", 
    x"447a", x"4478", x"4475", x"4472", x"4470", x"446d", x"446a", x"4468", 
    x"4465", x"4462", x"4460", x"445d", x"445a", x"4458", x"4455", x"4452", 
    x"4450", x"444d", x"444a", x"4448", x"4445", x"4442", x"4440", x"443d", 
    x"443b", x"4438", x"4435", x"4433", x"4430", x"442d", x"442b", x"4428", 
    x"4425", x"4423", x"4420", x"441d", x"441b", x"4418", x"4415", x"4413", 
    x"4410", x"440d", x"440b", x"4408", x"4405", x"4403", x"4400", x"43fd", 
    x"43fb", x"43f8", x"43f5", x"43f3", x"43f0", x"43ed", x"43eb", x"43e8", 
    x"43e5", x"43e3", x"43e0", x"43dd", x"43db", x"43d8", x"43d5", x"43d3", 
    x"43d0", x"43cd", x"43cb", x"43c8", x"43c5", x"43c3", x"43c0", x"43bd", 
    x"43bb", x"43b8", x"43b5", x"43b3", x"43b0", x"43ad", x"43ab", x"43a8", 
    x"43a5", x"43a3", x"43a0", x"439d", x"439b", x"4398", x"4395", x"4393", 
    x"4390", x"438d", x"438b", x"4388", x"4385", x"4383", x"4380", x"437d", 
    x"437b", x"4378", x"4375", x"4373", x"4370", x"436d", x"436b", x"4368", 
    x"4365", x"4363", x"4360", x"435d", x"435b", x"4358", x"4355", x"4353", 
    x"4350", x"434d", x"434b", x"4348", x"4345", x"4343", x"4340", x"433d", 
    x"433b", x"4338", x"4335", x"4333", x"4330", x"432d", x"432b", x"4328", 
    x"4325", x"4323", x"4320", x"431d", x"431b", x"4318", x"4315", x"4313", 
    x"4310", x"430d", x"430a", x"4308", x"4305", x"4302", x"4300", x"42fd", 
    x"42fa", x"42f8", x"42f5", x"42f2", x"42f0", x"42ed", x"42ea", x"42e8", 
    x"42e5", x"42e2", x"42e0", x"42dd", x"42da", x"42d8", x"42d5", x"42d2", 
    x"42d0", x"42cd", x"42ca", x"42c8", x"42c5", x"42c2", x"42bf", x"42bd", 
    x"42ba", x"42b7", x"42b5", x"42b2", x"42af", x"42ad", x"42aa", x"42a7", 
    x"42a5", x"42a2", x"429f", x"429d", x"429a", x"4297", x"4295", x"4292", 
    x"428f", x"428d", x"428a", x"4287", x"4284", x"4282", x"427f", x"427c", 
    x"427a", x"4277", x"4274", x"4272", x"426f", x"426c", x"426a", x"4267", 
    x"4264", x"4262", x"425f", x"425c", x"425a", x"4257", x"4254", x"4251", 
    x"424f", x"424c", x"4249", x"4247", x"4244", x"4241", x"423f", x"423c", 
    x"4239", x"4237", x"4234", x"4231", x"422f", x"422c", x"4229", x"4226", 
    x"4224", x"4221", x"421e", x"421c", x"4219", x"4216", x"4214", x"4211", 
    x"420e", x"420c", x"4209", x"4206", x"4203", x"4201", x"41fe", x"41fb", 
    x"41f9", x"41f6", x"41f3", x"41f1", x"41ee", x"41eb", x"41e9", x"41e6", 
    x"41e3", x"41e0", x"41de", x"41db", x"41d8", x"41d6", x"41d3", x"41d0", 
    x"41ce", x"41cb", x"41c8", x"41c6", x"41c3", x"41c0", x"41bd", x"41bb", 
    x"41b8", x"41b5", x"41b3", x"41b0", x"41ad", x"41ab", x"41a8", x"41a5", 
    x"41a2", x"41a0", x"419d", x"419a", x"4198", x"4195", x"4192", x"4190", 
    x"418d", x"418a", x"4187", x"4185", x"4182", x"417f", x"417d", x"417a", 
    x"4177", x"4175", x"4172", x"416f", x"416d", x"416a", x"4167", x"4164", 
    x"4162", x"415f", x"415c", x"415a", x"4157", x"4154", x"4151", x"414f", 
    x"414c", x"4149", x"4147", x"4144", x"4141", x"413f", x"413c", x"4139", 
    x"4136", x"4134", x"4131", x"412e", x"412c", x"4129", x"4126", x"4124", 
    x"4121", x"411e", x"411b", x"4119", x"4116", x"4113", x"4111", x"410e", 
    x"410b", x"4108", x"4106", x"4103", x"4100", x"40fe", x"40fb", x"40f8", 
    x"40f6", x"40f3", x"40f0", x"40ed", x"40eb", x"40e8", x"40e5", x"40e3", 
    x"40e0", x"40dd", x"40da", x"40d8", x"40d5", x"40d2", x"40d0", x"40cd", 
    x"40ca", x"40c8", x"40c5", x"40c2", x"40bf", x"40bd", x"40ba", x"40b7", 
    x"40b5", x"40b2", x"40af", x"40ac", x"40aa", x"40a7", x"40a4", x"40a2", 
    x"409f", x"409c", x"4099", x"4097", x"4094", x"4091", x"408f", x"408c", 
    x"4089", x"4086", x"4084", x"4081", x"407e", x"407c", x"4079", x"4076", 
    x"4073", x"4071", x"406e", x"406b", x"4069", x"4066", x"4063", x"4060", 
    x"405e", x"405b", x"4058", x"4056", x"4053", x"4050", x"404d", x"404b", 
    x"4048", x"4045", x"4043", x"4040", x"403d", x"403a", x"4038", x"4035", 
    x"4032", x"4030", x"402d", x"402a", x"4027", x"4025", x"4022", x"401f", 
    x"401d", x"401a", x"4017", x"4014", x"4012", x"400f", x"400c", x"4009", 
    x"4007", x"4004", x"4001", x"3fff", x"3ffc", x"3ff9", x"3ff6", x"3ff4", 
    x"3ff1", x"3fee", x"3fec", x"3fe9", x"3fe6", x"3fe3", x"3fe1", x"3fde", 
    x"3fdb", x"3fd8", x"3fd6", x"3fd3", x"3fd0", x"3fce", x"3fcb", x"3fc8", 
    x"3fc5", x"3fc3", x"3fc0", x"3fbd", x"3fbb", x"3fb8", x"3fb5", x"3fb2", 
    x"3fb0", x"3fad", x"3faa", x"3fa7", x"3fa5", x"3fa2", x"3f9f", x"3f9d", 
    x"3f9a", x"3f97", x"3f94", x"3f92", x"3f8f", x"3f8c", x"3f89", x"3f87", 
    x"3f84", x"3f81", x"3f7f", x"3f7c", x"3f79", x"3f76", x"3f74", x"3f71", 
    x"3f6e", x"3f6b", x"3f69", x"3f66", x"3f63", x"3f61", x"3f5e", x"3f5b", 
    x"3f58", x"3f56", x"3f53", x"3f50", x"3f4d", x"3f4b", x"3f48", x"3f45", 
    x"3f43", x"3f40", x"3f3d", x"3f3a", x"3f38", x"3f35", x"3f32", x"3f2f", 
    x"3f2d", x"3f2a", x"3f27", x"3f24", x"3f22", x"3f1f", x"3f1c", x"3f1a", 
    x"3f17", x"3f14", x"3f11", x"3f0f", x"3f0c", x"3f09", x"3f06", x"3f04", 
    x"3f01", x"3efe", x"3efb", x"3ef9", x"3ef6", x"3ef3", x"3ef1", x"3eee", 
    x"3eeb", x"3ee8", x"3ee6", x"3ee3", x"3ee0", x"3edd", x"3edb", x"3ed8", 
    x"3ed5", x"3ed2", x"3ed0", x"3ecd", x"3eca", x"3ec7", x"3ec5", x"3ec2", 
    x"3ebf", x"3ebd", x"3eba", x"3eb7", x"3eb4", x"3eb2", x"3eaf", x"3eac", 
    x"3ea9", x"3ea7", x"3ea4", x"3ea1", x"3e9e", x"3e9c", x"3e99", x"3e96", 
    x"3e93", x"3e91", x"3e8e", x"3e8b", x"3e88", x"3e86", x"3e83", x"3e80", 
    x"3e7d", x"3e7b", x"3e78", x"3e75", x"3e73", x"3e70", x"3e6d", x"3e6a", 
    x"3e68", x"3e65", x"3e62", x"3e5f", x"3e5d", x"3e5a", x"3e57", x"3e54", 
    x"3e52", x"3e4f", x"3e4c", x"3e49", x"3e47", x"3e44", x"3e41", x"3e3e", 
    x"3e3c", x"3e39", x"3e36", x"3e33", x"3e31", x"3e2e", x"3e2b", x"3e28", 
    x"3e26", x"3e23", x"3e20", x"3e1d", x"3e1b", x"3e18", x"3e15", x"3e12", 
    x"3e10", x"3e0d", x"3e0a", x"3e07", x"3e05", x"3e02", x"3dff", x"3dfc", 
    x"3dfa", x"3df7", x"3df4", x"3df1", x"3def", x"3dec", x"3de9", x"3de6", 
    x"3de4", x"3de1", x"3dde", x"3ddb", x"3dd9", x"3dd6", x"3dd3", x"3dd0", 
    x"3dce", x"3dcb", x"3dc8", x"3dc5", x"3dc3", x"3dc0", x"3dbd", x"3dba", 
    x"3db8", x"3db5", x"3db2", x"3daf", x"3dad", x"3daa", x"3da7", x"3da4", 
    x"3da2", x"3d9f", x"3d9c", x"3d99", x"3d97", x"3d94", x"3d91", x"3d8e", 
    x"3d8c", x"3d89", x"3d86", x"3d83", x"3d81", x"3d7e", x"3d7b", x"3d78", 
    x"3d76", x"3d73", x"3d70", x"3d6d", x"3d6b", x"3d68", x"3d65", x"3d62", 
    x"3d60", x"3d5d", x"3d5a", x"3d57", x"3d55", x"3d52", x"3d4f", x"3d4c", 
    x"3d4a", x"3d47", x"3d44", x"3d41", x"3d3e", x"3d3c", x"3d39", x"3d36", 
    x"3d33", x"3d31", x"3d2e", x"3d2b", x"3d28", x"3d26", x"3d23", x"3d20", 
    x"3d1d", x"3d1b", x"3d18", x"3d15", x"3d12", x"3d10", x"3d0d", x"3d0a", 
    x"3d07", x"3d05", x"3d02", x"3cff", x"3cfc", x"3cf9", x"3cf7", x"3cf4", 
    x"3cf1", x"3cee", x"3cec", x"3ce9", x"3ce6", x"3ce3", x"3ce1", x"3cde", 
    x"3cdb", x"3cd8", x"3cd6", x"3cd3", x"3cd0", x"3ccd", x"3cca", x"3cc8", 
    x"3cc5", x"3cc2", x"3cbf", x"3cbd", x"3cba", x"3cb7", x"3cb4", x"3cb2", 
    x"3caf", x"3cac", x"3ca9", x"3ca7", x"3ca4", x"3ca1", x"3c9e", x"3c9b", 
    x"3c99", x"3c96", x"3c93", x"3c90", x"3c8e", x"3c8b", x"3c88", x"3c85", 
    x"3c83", x"3c80", x"3c7d", x"3c7a", x"3c77", x"3c75", x"3c72", x"3c6f", 
    x"3c6c", x"3c6a", x"3c67", x"3c64", x"3c61", x"3c5f", x"3c5c", x"3c59", 
    x"3c56", x"3c53", x"3c51", x"3c4e", x"3c4b", x"3c48", x"3c46", x"3c43", 
    x"3c40", x"3c3d", x"3c3b", x"3c38", x"3c35", x"3c32", x"3c2f", x"3c2d", 
    x"3c2a", x"3c27", x"3c24", x"3c22", x"3c1f", x"3c1c", x"3c19", x"3c16", 
    x"3c14", x"3c11", x"3c0e", x"3c0b", x"3c09", x"3c06", x"3c03", x"3c00", 
    x"3bfe", x"3bfb", x"3bf8", x"3bf5", x"3bf2", x"3bf0", x"3bed", x"3bea", 
    x"3be7", x"3be5", x"3be2", x"3bdf", x"3bdc", x"3bd9", x"3bd7", x"3bd4", 
    x"3bd1", x"3bce", x"3bcc", x"3bc9", x"3bc6", x"3bc3", x"3bc0", x"3bbe", 
    x"3bbb", x"3bb8", x"3bb5", x"3bb3", x"3bb0", x"3bad", x"3baa", x"3ba7", 
    x"3ba5", x"3ba2", x"3b9f", x"3b9c", x"3b9a", x"3b97", x"3b94", x"3b91", 
    x"3b8e", x"3b8c", x"3b89", x"3b86", x"3b83", x"3b81", x"3b7e", x"3b7b", 
    x"3b78", x"3b75", x"3b73", x"3b70", x"3b6d", x"3b6a", x"3b67", x"3b65", 
    x"3b62", x"3b5f", x"3b5c", x"3b5a", x"3b57", x"3b54", x"3b51", x"3b4e", 
    x"3b4c", x"3b49", x"3b46", x"3b43", x"3b40", x"3b3e", x"3b3b", x"3b38", 
    x"3b35", x"3b33", x"3b30", x"3b2d", x"3b2a", x"3b27", x"3b25", x"3b22", 
    x"3b1f", x"3b1c", x"3b19", x"3b17", x"3b14", x"3b11", x"3b0e", x"3b0c", 
    x"3b09", x"3b06", x"3b03", x"3b00", x"3afe", x"3afb", x"3af8", x"3af5", 
    x"3af2", x"3af0", x"3aed", x"3aea", x"3ae7", x"3ae5", x"3ae2", x"3adf", 
    x"3adc", x"3ad9", x"3ad7", x"3ad4", x"3ad1", x"3ace", x"3acb", x"3ac9", 
    x"3ac6", x"3ac3", x"3ac0", x"3abd", x"3abb", x"3ab8", x"3ab5", x"3ab2", 
    x"3ab0", x"3aad", x"3aaa", x"3aa7", x"3aa4", x"3aa2", x"3a9f", x"3a9c", 
    x"3a99", x"3a96", x"3a94", x"3a91", x"3a8e", x"3a8b", x"3a88", x"3a86", 
    x"3a83", x"3a80", x"3a7d", x"3a7a", x"3a78", x"3a75", x"3a72", x"3a6f", 
    x"3a6c", x"3a6a", x"3a67", x"3a64", x"3a61", x"3a5e", x"3a5c", x"3a59", 
    x"3a56", x"3a53", x"3a51", x"3a4e", x"3a4b", x"3a48", x"3a45", x"3a43", 
    x"3a40", x"3a3d", x"3a3a", x"3a37", x"3a35", x"3a32", x"3a2f", x"3a2c", 
    x"3a29", x"3a27", x"3a24", x"3a21", x"3a1e", x"3a1b", x"3a19", x"3a16", 
    x"3a13", x"3a10", x"3a0d", x"3a0b", x"3a08", x"3a05", x"3a02", x"39ff", 
    x"39fd", x"39fa", x"39f7", x"39f4", x"39f1", x"39ef", x"39ec", x"39e9", 
    x"39e6", x"39e3", x"39e1", x"39de", x"39db", x"39d8", x"39d5", x"39d3", 
    x"39d0", x"39cd", x"39ca", x"39c7", x"39c5", x"39c2", x"39bf", x"39bc", 
    x"39b9", x"39b6", x"39b4", x"39b1", x"39ae", x"39ab", x"39a8", x"39a6", 
    x"39a3", x"39a0", x"399d", x"399a", x"3998", x"3995", x"3992", x"398f", 
    x"398c", x"398a", x"3987", x"3984", x"3981", x"397e", x"397c", x"3979", 
    x"3976", x"3973", x"3970", x"396e", x"396b", x"3968", x"3965", x"3962", 
    x"3960", x"395d", x"395a", x"3957", x"3954", x"3951", x"394f", x"394c", 
    x"3949", x"3946", x"3943", x"3941", x"393e", x"393b", x"3938", x"3935", 
    x"3933", x"3930", x"392d", x"392a", x"3927", x"3924", x"3922", x"391f", 
    x"391c", x"3919", x"3916", x"3914", x"3911", x"390e", x"390b", x"3908", 
    x"3906", x"3903", x"3900", x"38fd", x"38fa", x"38f8", x"38f5", x"38f2", 
    x"38ef", x"38ec", x"38e9", x"38e7", x"38e4", x"38e1", x"38de", x"38db", 
    x"38d9", x"38d6", x"38d3", x"38d0", x"38cd", x"38ca", x"38c8", x"38c5", 
    x"38c2", x"38bf", x"38bc", x"38ba", x"38b7", x"38b4", x"38b1", x"38ae", 
    x"38ab", x"38a9", x"38a6", x"38a3", x"38a0", x"389d", x"389b", x"3898", 
    x"3895", x"3892", x"388f", x"388d", x"388a", x"3887", x"3884", x"3881", 
    x"387e", x"387c", x"3879", x"3876", x"3873", x"3870", x"386d", x"386b", 
    x"3868", x"3865", x"3862", x"385f", x"385d", x"385a", x"3857", x"3854", 
    x"3851", x"384e", x"384c", x"3849", x"3846", x"3843", x"3840", x"383e", 
    x"383b", x"3838", x"3835", x"3832", x"382f", x"382d", x"382a", x"3827", 
    x"3824", x"3821", x"381e", x"381c", x"3819", x"3816", x"3813", x"3810", 
    x"380e", x"380b", x"3808", x"3805", x"3802", x"37ff", x"37fd", x"37fa", 
    x"37f7", x"37f4", x"37f1", x"37ee", x"37ec", x"37e9", x"37e6", x"37e3", 
    x"37e0", x"37de", x"37db", x"37d8", x"37d5", x"37d2", x"37cf", x"37cd", 
    x"37ca", x"37c7", x"37c4", x"37c1", x"37be", x"37bc", x"37b9", x"37b6", 
    x"37b3", x"37b0", x"37ad", x"37ab", x"37a8", x"37a5", x"37a2", x"379f", 
    x"379c", x"379a", x"3797", x"3794", x"3791", x"378e", x"378b", x"3789", 
    x"3786", x"3783", x"3780", x"377d", x"377b", x"3778", x"3775", x"3772", 
    x"376f", x"376c", x"376a", x"3767", x"3764", x"3761", x"375e", x"375b", 
    x"3759", x"3756", x"3753", x"3750", x"374d", x"374a", x"3748", x"3745", 
    x"3742", x"373f", x"373c", x"3739", x"3737", x"3734", x"3731", x"372e", 
    x"372b", x"3728", x"3726", x"3723", x"3720", x"371d", x"371a", x"3717", 
    x"3715", x"3712", x"370f", x"370c", x"3709", x"3706", x"3703", x"3701", 
    x"36fe", x"36fb", x"36f8", x"36f5", x"36f2", x"36f0", x"36ed", x"36ea", 
    x"36e7", x"36e4", x"36e1", x"36df", x"36dc", x"36d9", x"36d6", x"36d3", 
    x"36d0", x"36ce", x"36cb", x"36c8", x"36c5", x"36c2", x"36bf", x"36bd", 
    x"36ba", x"36b7", x"36b4", x"36b1", x"36ae", x"36ab", x"36a9", x"36a6", 
    x"36a3", x"36a0", x"369d", x"369a", x"3698", x"3695", x"3692", x"368f", 
    x"368c", x"3689", x"3687", x"3684", x"3681", x"367e", x"367b", x"3678", 
    x"3676", x"3673", x"3670", x"366d", x"366a", x"3667", x"3664", x"3662", 
    x"365f", x"365c", x"3659", x"3656", x"3653", x"3651", x"364e", x"364b", 
    x"3648", x"3645", x"3642", x"363f", x"363d", x"363a", x"3637", x"3634", 
    x"3631", x"362e", x"362c", x"3629", x"3626", x"3623", x"3620", x"361d", 
    x"361a", x"3618", x"3615", x"3612", x"360f", x"360c", x"3609", x"3607", 
    x"3604", x"3601", x"35fe", x"35fb", x"35f8", x"35f5", x"35f3", x"35f0", 
    x"35ed", x"35ea", x"35e7", x"35e4", x"35e1", x"35df", x"35dc", x"35d9", 
    x"35d6", x"35d3", x"35d0", x"35ce", x"35cb", x"35c8", x"35c5", x"35c2", 
    x"35bf", x"35bc", x"35ba", x"35b7", x"35b4", x"35b1", x"35ae", x"35ab", 
    x"35a8", x"35a6", x"35a3", x"35a0", x"359d", x"359a", x"3597", x"3595", 
    x"3592", x"358f", x"358c", x"3589", x"3586", x"3583", x"3581", x"357e", 
    x"357b", x"3578", x"3575", x"3572", x"356f", x"356d", x"356a", x"3567", 
    x"3564", x"3561", x"355e", x"355b", x"3559", x"3556", x"3553", x"3550", 
    x"354d", x"354a", x"3547", x"3545", x"3542", x"353f", x"353c", x"3539", 
    x"3536", x"3533", x"3531", x"352e", x"352b", x"3528", x"3525", x"3522", 
    x"351f", x"351d", x"351a", x"3517", x"3514", x"3511", x"350e", x"350b", 
    x"3509", x"3506", x"3503", x"3500", x"34fd", x"34fa", x"34f7", x"34f5", 
    x"34f2", x"34ef", x"34ec", x"34e9", x"34e6", x"34e3", x"34e1", x"34de", 
    x"34db", x"34d8", x"34d5", x"34d2", x"34cf", x"34cc", x"34ca", x"34c7", 
    x"34c4", x"34c1", x"34be", x"34bb", x"34b8", x"34b6", x"34b3", x"34b0", 
    x"34ad", x"34aa", x"34a7", x"34a4", x"34a2", x"349f", x"349c", x"3499", 
    x"3496", x"3493", x"3490", x"348e", x"348b", x"3488", x"3485", x"3482", 
    x"347f", x"347c", x"3479", x"3477", x"3474", x"3471", x"346e", x"346b", 
    x"3468", x"3465", x"3463", x"3460", x"345d", x"345a", x"3457", x"3454", 
    x"3451", x"344e", x"344c", x"3449", x"3446", x"3443", x"3440", x"343d", 
    x"343a", x"3438", x"3435", x"3432", x"342f", x"342c", x"3429", x"3426", 
    x"3423", x"3421", x"341e", x"341b", x"3418", x"3415", x"3412", x"340f", 
    x"340c", x"340a", x"3407", x"3404", x"3401", x"33fe", x"33fb", x"33f8", 
    x"33f6", x"33f3", x"33f0", x"33ed", x"33ea", x"33e7", x"33e4", x"33e1", 
    x"33df", x"33dc", x"33d9", x"33d6", x"33d3", x"33d0", x"33cd", x"33ca", 
    x"33c8", x"33c5", x"33c2", x"33bf", x"33bc", x"33b9", x"33b6", x"33b3", 
    x"33b1", x"33ae", x"33ab", x"33a8", x"33a5", x"33a2", x"339f", x"339c", 
    x"339a", x"3397", x"3394", x"3391", x"338e", x"338b", x"3388", x"3385", 
    x"3383", x"3380", x"337d", x"337a", x"3377", x"3374", x"3371", x"336e", 
    x"336c", x"3369", x"3366", x"3363", x"3360", x"335d", x"335a", x"3357", 
    x"3355", x"3352", x"334f", x"334c", x"3349", x"3346", x"3343", x"3340", 
    x"333e", x"333b", x"3338", x"3335", x"3332", x"332f", x"332c", x"3329", 
    x"3326", x"3324", x"3321", x"331e", x"331b", x"3318", x"3315", x"3312", 
    x"330f", x"330d", x"330a", x"3307", x"3304", x"3301", x"32fe", x"32fb", 
    x"32f8", x"32f6", x"32f3", x"32f0", x"32ed", x"32ea", x"32e7", x"32e4", 
    x"32e1", x"32de", x"32dc", x"32d9", x"32d6", x"32d3", x"32d0", x"32cd", 
    x"32ca", x"32c7", x"32c5", x"32c2", x"32bf", x"32bc", x"32b9", x"32b6", 
    x"32b3", x"32b0", x"32ad", x"32ab", x"32a8", x"32a5", x"32a2", x"329f", 
    x"329c", x"3299", x"3296", x"3293", x"3291", x"328e", x"328b", x"3288", 
    x"3285", x"3282", x"327f", x"327c", x"3279", x"3277", x"3274", x"3271", 
    x"326e", x"326b", x"3268", x"3265", x"3262", x"325f", x"325d", x"325a", 
    x"3257", x"3254", x"3251", x"324e", x"324b", x"3248", x"3246", x"3243", 
    x"3240", x"323d", x"323a", x"3237", x"3234", x"3231", x"322e", x"322b", 
    x"3229", x"3226", x"3223", x"3220", x"321d", x"321a", x"3217", x"3214", 
    x"3211", x"320f", x"320c", x"3209", x"3206", x"3203", x"3200", x"31fd", 
    x"31fa", x"31f7", x"31f5", x"31f2", x"31ef", x"31ec", x"31e9", x"31e6", 
    x"31e3", x"31e0", x"31dd", x"31db", x"31d8", x"31d5", x"31d2", x"31cf", 
    x"31cc", x"31c9", x"31c6", x"31c3", x"31c0", x"31be", x"31bb", x"31b8", 
    x"31b5", x"31b2", x"31af", x"31ac", x"31a9", x"31a6", x"31a4", x"31a1", 
    x"319e", x"319b", x"3198", x"3195", x"3192", x"318f", x"318c", x"3189", 
    x"3187", x"3184", x"3181", x"317e", x"317b", x"3178", x"3175", x"3172", 
    x"316f", x"316c", x"316a", x"3167", x"3164", x"3161", x"315e", x"315b", 
    x"3158", x"3155", x"3152", x"3150", x"314d", x"314a", x"3147", x"3144", 
    x"3141", x"313e", x"313b", x"3138", x"3135", x"3133", x"3130", x"312d", 
    x"312a", x"3127", x"3124", x"3121", x"311e", x"311b", x"3118", x"3116", 
    x"3113", x"3110", x"310d", x"310a", x"3107", x"3104", x"3101", x"30fe", 
    x"30fb", x"30f8", x"30f6", x"30f3", x"30f0", x"30ed", x"30ea", x"30e7", 
    x"30e4", x"30e1", x"30de", x"30db", x"30d9", x"30d6", x"30d3", x"30d0", 
    x"30cd", x"30ca", x"30c7", x"30c4", x"30c1", x"30be", x"30bc", x"30b9", 
    x"30b6", x"30b3", x"30b0", x"30ad", x"30aa", x"30a7", x"30a4", x"30a1", 
    x"309e", x"309c", x"3099", x"3096", x"3093", x"3090", x"308d", x"308a", 
    x"3087", x"3084", x"3081", x"307e", x"307c", x"3079", x"3076", x"3073", 
    x"3070", x"306d", x"306a", x"3067", x"3064", x"3061", x"305e", x"305c", 
    x"3059", x"3056", x"3053", x"3050", x"304d", x"304a", x"3047", x"3044", 
    x"3041", x"303e", x"303c", x"3039", x"3036", x"3033", x"3030", x"302d", 
    x"302a", x"3027", x"3024", x"3021", x"301e", x"301c", x"3019", x"3016", 
    x"3013", x"3010", x"300d", x"300a", x"3007", x"3004", x"3001", x"2ffe", 
    x"2ffc", x"2ff9", x"2ff6", x"2ff3", x"2ff0", x"2fed", x"2fea", x"2fe7", 
    x"2fe4", x"2fe1", x"2fde", x"2fdb", x"2fd9", x"2fd6", x"2fd3", x"2fd0", 
    x"2fcd", x"2fca", x"2fc7", x"2fc4", x"2fc1", x"2fbe", x"2fbb", x"2fb9", 
    x"2fb6", x"2fb3", x"2fb0", x"2fad", x"2faa", x"2fa7", x"2fa4", x"2fa1", 
    x"2f9e", x"2f9b", x"2f98", x"2f96", x"2f93", x"2f90", x"2f8d", x"2f8a", 
    x"2f87", x"2f84", x"2f81", x"2f7e", x"2f7b", x"2f78", x"2f75", x"2f73", 
    x"2f70", x"2f6d", x"2f6a", x"2f67", x"2f64", x"2f61", x"2f5e", x"2f5b", 
    x"2f58", x"2f55", x"2f52", x"2f50", x"2f4d", x"2f4a", x"2f47", x"2f44", 
    x"2f41", x"2f3e", x"2f3b", x"2f38", x"2f35", x"2f32", x"2f2f", x"2f2c", 
    x"2f2a", x"2f27", x"2f24", x"2f21", x"2f1e", x"2f1b", x"2f18", x"2f15", 
    x"2f12", x"2f0f", x"2f0c", x"2f09", x"2f06", x"2f04", x"2f01", x"2efe", 
    x"2efb", x"2ef8", x"2ef5", x"2ef2", x"2eef", x"2eec", x"2ee9", x"2ee6", 
    x"2ee3", x"2ee1", x"2ede", x"2edb", x"2ed8", x"2ed5", x"2ed2", x"2ecf", 
    x"2ecc", x"2ec9", x"2ec6", x"2ec3", x"2ec0", x"2ebd", x"2eba", x"2eb8", 
    x"2eb5", x"2eb2", x"2eaf", x"2eac", x"2ea9", x"2ea6", x"2ea3", x"2ea0", 
    x"2e9d", x"2e9a", x"2e97", x"2e94", x"2e92", x"2e8f", x"2e8c", x"2e89", 
    x"2e86", x"2e83", x"2e80", x"2e7d", x"2e7a", x"2e77", x"2e74", x"2e71", 
    x"2e6e", x"2e6b", x"2e69", x"2e66", x"2e63", x"2e60", x"2e5d", x"2e5a", 
    x"2e57", x"2e54", x"2e51", x"2e4e", x"2e4b", x"2e48", x"2e45", x"2e42", 
    x"2e40", x"2e3d", x"2e3a", x"2e37", x"2e34", x"2e31", x"2e2e", x"2e2b", 
    x"2e28", x"2e25", x"2e22", x"2e1f", x"2e1c", x"2e19", x"2e17", x"2e14", 
    x"2e11", x"2e0e", x"2e0b", x"2e08", x"2e05", x"2e02", x"2dff", x"2dfc", 
    x"2df9", x"2df6", x"2df3", x"2df0", x"2dee", x"2deb", x"2de8", x"2de5", 
    x"2de2", x"2ddf", x"2ddc", x"2dd9", x"2dd6", x"2dd3", x"2dd0", x"2dcd", 
    x"2dca", x"2dc7", x"2dc4", x"2dc2", x"2dbf", x"2dbc", x"2db9", x"2db6", 
    x"2db3", x"2db0", x"2dad", x"2daa", x"2da7", x"2da4", x"2da1", x"2d9e", 
    x"2d9b", x"2d98", x"2d95", x"2d93", x"2d90", x"2d8d", x"2d8a", x"2d87", 
    x"2d84", x"2d81", x"2d7e", x"2d7b", x"2d78", x"2d75", x"2d72", x"2d6f", 
    x"2d6c", x"2d69", x"2d67", x"2d64", x"2d61", x"2d5e", x"2d5b", x"2d58", 
    x"2d55", x"2d52", x"2d4f", x"2d4c", x"2d49", x"2d46", x"2d43", x"2d40", 
    x"2d3d", x"2d3a", x"2d37", x"2d35", x"2d32", x"2d2f", x"2d2c", x"2d29", 
    x"2d26", x"2d23", x"2d20", x"2d1d", x"2d1a", x"2d17", x"2d14", x"2d11", 
    x"2d0e", x"2d0b", x"2d08", x"2d06", x"2d03", x"2d00", x"2cfd", x"2cfa", 
    x"2cf7", x"2cf4", x"2cf1", x"2cee", x"2ceb", x"2ce8", x"2ce5", x"2ce2", 
    x"2cdf", x"2cdc", x"2cd9", x"2cd6", x"2cd4", x"2cd1", x"2cce", x"2ccb", 
    x"2cc8", x"2cc5", x"2cc2", x"2cbf", x"2cbc", x"2cb9", x"2cb6", x"2cb3", 
    x"2cb0", x"2cad", x"2caa", x"2ca7", x"2ca4", x"2ca1", x"2c9f", x"2c9c", 
    x"2c99", x"2c96", x"2c93", x"2c90", x"2c8d", x"2c8a", x"2c87", x"2c84", 
    x"2c81", x"2c7e", x"2c7b", x"2c78", x"2c75", x"2c72", x"2c6f", x"2c6c", 
    x"2c6a", x"2c67", x"2c64", x"2c61", x"2c5e", x"2c5b", x"2c58", x"2c55", 
    x"2c52", x"2c4f", x"2c4c", x"2c49", x"2c46", x"2c43", x"2c40", x"2c3d", 
    x"2c3a", x"2c37", x"2c34", x"2c32", x"2c2f", x"2c2c", x"2c29", x"2c26", 
    x"2c23", x"2c20", x"2c1d", x"2c1a", x"2c17", x"2c14", x"2c11", x"2c0e", 
    x"2c0b", x"2c08", x"2c05", x"2c02", x"2bff", x"2bfc", x"2bf9", x"2bf7", 
    x"2bf4", x"2bf1", x"2bee", x"2beb", x"2be8", x"2be5", x"2be2", x"2bdf", 
    x"2bdc", x"2bd9", x"2bd6", x"2bd3", x"2bd0", x"2bcd", x"2bca", x"2bc7", 
    x"2bc4", x"2bc1", x"2bbe", x"2bbb", x"2bb9", x"2bb6", x"2bb3", x"2bb0", 
    x"2bad", x"2baa", x"2ba7", x"2ba4", x"2ba1", x"2b9e", x"2b9b", x"2b98", 
    x"2b95", x"2b92", x"2b8f", x"2b8c", x"2b89", x"2b86", x"2b83", x"2b80", 
    x"2b7d", x"2b7b", x"2b78", x"2b75", x"2b72", x"2b6f", x"2b6c", x"2b69", 
    x"2b66", x"2b63", x"2b60", x"2b5d", x"2b5a", x"2b57", x"2b54", x"2b51", 
    x"2b4e", x"2b4b", x"2b48", x"2b45", x"2b42", x"2b3f", x"2b3c", x"2b39", 
    x"2b37", x"2b34", x"2b31", x"2b2e", x"2b2b", x"2b28", x"2b25", x"2b22", 
    x"2b1f", x"2b1c", x"2b19", x"2b16", x"2b13", x"2b10", x"2b0d", x"2b0a", 
    x"2b07", x"2b04", x"2b01", x"2afe", x"2afb", x"2af8", x"2af5", x"2af2", 
    x"2af0", x"2aed", x"2aea", x"2ae7", x"2ae4", x"2ae1", x"2ade", x"2adb", 
    x"2ad8", x"2ad5", x"2ad2", x"2acf", x"2acc", x"2ac9", x"2ac6", x"2ac3", 
    x"2ac0", x"2abd", x"2aba", x"2ab7", x"2ab4", x"2ab1", x"2aae", x"2aab", 
    x"2aa8", x"2aa6", x"2aa3", x"2aa0", x"2a9d", x"2a9a", x"2a97", x"2a94", 
    x"2a91", x"2a8e", x"2a8b", x"2a88", x"2a85", x"2a82", x"2a7f", x"2a7c", 
    x"2a79", x"2a76", x"2a73", x"2a70", x"2a6d", x"2a6a", x"2a67", x"2a64", 
    x"2a61", x"2a5e", x"2a5b", x"2a58", x"2a56", x"2a53", x"2a50", x"2a4d", 
    x"2a4a", x"2a47", x"2a44", x"2a41", x"2a3e", x"2a3b", x"2a38", x"2a35", 
    x"2a32", x"2a2f", x"2a2c", x"2a29", x"2a26", x"2a23", x"2a20", x"2a1d", 
    x"2a1a", x"2a17", x"2a14", x"2a11", x"2a0e", x"2a0b", x"2a08", x"2a05", 
    x"2a02", x"29ff", x"29fd", x"29fa", x"29f7", x"29f4", x"29f1", x"29ee", 
    x"29eb", x"29e8", x"29e5", x"29e2", x"29df", x"29dc", x"29d9", x"29d6", 
    x"29d3", x"29d0", x"29cd", x"29ca", x"29c7", x"29c4", x"29c1", x"29be", 
    x"29bb", x"29b8", x"29b5", x"29b2", x"29af", x"29ac", x"29a9", x"29a6", 
    x"29a3", x"29a0", x"299e", x"299b", x"2998", x"2995", x"2992", x"298f", 
    x"298c", x"2989", x"2986", x"2983", x"2980", x"297d", x"297a", x"2977", 
    x"2974", x"2971", x"296e", x"296b", x"2968", x"2965", x"2962", x"295f", 
    x"295c", x"2959", x"2956", x"2953", x"2950", x"294d", x"294a", x"2947", 
    x"2944", x"2941", x"293e", x"293b", x"2938", x"2935", x"2932", x"2930", 
    x"292d", x"292a", x"2927", x"2924", x"2921", x"291e", x"291b", x"2918", 
    x"2915", x"2912", x"290f", x"290c", x"2909", x"2906", x"2903", x"2900", 
    x"28fd", x"28fa", x"28f7", x"28f4", x"28f1", x"28ee", x"28eb", x"28e8", 
    x"28e5", x"28e2", x"28df", x"28dc", x"28d9", x"28d6", x"28d3", x"28d0", 
    x"28cd", x"28ca", x"28c7", x"28c4", x"28c1", x"28be", x"28bb", x"28b8", 
    x"28b5", x"28b3", x"28b0", x"28ad", x"28aa", x"28a7", x"28a4", x"28a1", 
    x"289e", x"289b", x"2898", x"2895", x"2892", x"288f", x"288c", x"2889", 
    x"2886", x"2883", x"2880", x"287d", x"287a", x"2877", x"2874", x"2871", 
    x"286e", x"286b", x"2868", x"2865", x"2862", x"285f", x"285c", x"2859", 
    x"2856", x"2853", x"2850", x"284d", x"284a", x"2847", x"2844", x"2841", 
    x"283e", x"283b", x"2838", x"2835", x"2832", x"282f", x"282c", x"2829", 
    x"2826", x"2823", x"2820", x"281d", x"281a", x"2817", x"2815", x"2812", 
    x"280f", x"280c", x"2809", x"2806", x"2803", x"2800", x"27fd", x"27fa", 
    x"27f7", x"27f4", x"27f1", x"27ee", x"27eb", x"27e8", x"27e5", x"27e2", 
    x"27df", x"27dc", x"27d9", x"27d6", x"27d3", x"27d0", x"27cd", x"27ca", 
    x"27c7", x"27c4", x"27c1", x"27be", x"27bb", x"27b8", x"27b5", x"27b2", 
    x"27af", x"27ac", x"27a9", x"27a6", x"27a3", x"27a0", x"279d", x"279a", 
    x"2797", x"2794", x"2791", x"278e", x"278b", x"2788", x"2785", x"2782", 
    x"277f", x"277c", x"2779", x"2776", x"2773", x"2770", x"276d", x"276a", 
    x"2767", x"2764", x"2761", x"275e", x"275b", x"2758", x"2755", x"2752", 
    x"274f", x"274c", x"2749", x"2746", x"2743", x"2740", x"273d", x"273a", 
    x"2737", x"2734", x"2731", x"272f", x"272c", x"2729", x"2726", x"2723", 
    x"2720", x"271d", x"271a", x"2717", x"2714", x"2711", x"270e", x"270b", 
    x"2708", x"2705", x"2702", x"26ff", x"26fc", x"26f9", x"26f6", x"26f3", 
    x"26f0", x"26ed", x"26ea", x"26e7", x"26e4", x"26e1", x"26de", x"26db", 
    x"26d8", x"26d5", x"26d2", x"26cf", x"26cc", x"26c9", x"26c6", x"26c3", 
    x"26c0", x"26bd", x"26ba", x"26b7", x"26b4", x"26b1", x"26ae", x"26ab", 
    x"26a8", x"26a5", x"26a2", x"269f", x"269c", x"2699", x"2696", x"2693", 
    x"2690", x"268d", x"268a", x"2687", x"2684", x"2681", x"267e", x"267b", 
    x"2678", x"2675", x"2672", x"266f", x"266c", x"2669", x"2666", x"2663", 
    x"2660", x"265d", x"265a", x"2657", x"2654", x"2651", x"264e", x"264b", 
    x"2648", x"2645", x"2642", x"263f", x"263c", x"2639", x"2636", x"2633", 
    x"2630", x"262d", x"262a", x"2627", x"2624", x"2621", x"261e", x"261b", 
    x"2618", x"2615", x"2612", x"260f", x"260c", x"2609", x"2606", x"2603", 
    x"2600", x"25fd", x"25fa", x"25f7", x"25f4", x"25f1", x"25ee", x"25eb", 
    x"25e8", x"25e5", x"25e2", x"25df", x"25dc", x"25d9", x"25d6", x"25d3", 
    x"25d0", x"25cd", x"25ca", x"25c7", x"25c4", x"25c1", x"25be", x"25bb", 
    x"25b8", x"25b5", x"25b2", x"25af", x"25ac", x"25a9", x"25a6", x"25a3", 
    x"25a0", x"259d", x"259a", x"2597", x"2594", x"2591", x"258e", x"258b", 
    x"2588", x"2585", x"2582", x"257f", x"257c", x"2579", x"2576", x"2573", 
    x"2570", x"256d", x"256a", x"2567", x"2564", x"2561", x"255e", x"255b", 
    x"2558", x"2555", x"2552", x"254f", x"254c", x"2549", x"2546", x"2543", 
    x"2540", x"253d", x"253a", x"2537", x"2534", x"2531", x"252e", x"252b", 
    x"2528", x"2525", x"2522", x"251f", x"251c", x"2519", x"2516", x"2513", 
    x"2510", x"250d", x"250a", x"2507", x"2504", x"2501", x"24fe", x"24fb", 
    x"24f8", x"24f5", x"24f2", x"24ef", x"24ec", x"24e9", x"24e6", x"24e3", 
    x"24e0", x"24dd", x"24da", x"24d7", x"24d4", x"24d1", x"24ce", x"24cb", 
    x"24c8", x"24c5", x"24c1", x"24be", x"24bb", x"24b8", x"24b5", x"24b2", 
    x"24af", x"24ac", x"24a9", x"24a6", x"24a3", x"24a0", x"249d", x"249a", 
    x"2497", x"2494", x"2491", x"248e", x"248b", x"2488", x"2485", x"2482", 
    x"247f", x"247c", x"2479", x"2476", x"2473", x"2470", x"246d", x"246a", 
    x"2467", x"2464", x"2461", x"245e", x"245b", x"2458", x"2455", x"2452", 
    x"244f", x"244c", x"2449", x"2446", x"2443", x"2440", x"243d", x"243a", 
    x"2437", x"2434", x"2431", x"242e", x"242b", x"2428", x"2425", x"2422", 
    x"241f", x"241c", x"2419", x"2416", x"2413", x"2410", x"240d", x"240a", 
    x"2407", x"2404", x"2401", x"23fe", x"23fb", x"23f8", x"23f5", x"23f2", 
    x"23ef", x"23ec", x"23e9", x"23e6", x"23e3", x"23e0", x"23dd", x"23da", 
    x"23d7", x"23d4", x"23d0", x"23cd", x"23ca", x"23c7", x"23c4", x"23c1", 
    x"23be", x"23bb", x"23b8", x"23b5", x"23b2", x"23af", x"23ac", x"23a9", 
    x"23a6", x"23a3", x"23a0", x"239d", x"239a", x"2397", x"2394", x"2391", 
    x"238e", x"238b", x"2388", x"2385", x"2382", x"237f", x"237c", x"2379", 
    x"2376", x"2373", x"2370", x"236d", x"236a", x"2367", x"2364", x"2361", 
    x"235e", x"235b", x"2358", x"2355", x"2352", x"234f", x"234c", x"2349", 
    x"2346", x"2343", x"2340", x"233d", x"233a", x"2337", x"2334", x"2331", 
    x"232e", x"232a", x"2327", x"2324", x"2321", x"231e", x"231b", x"2318", 
    x"2315", x"2312", x"230f", x"230c", x"2309", x"2306", x"2303", x"2300", 
    x"22fd", x"22fa", x"22f7", x"22f4", x"22f1", x"22ee", x"22eb", x"22e8", 
    x"22e5", x"22e2", x"22df", x"22dc", x"22d9", x"22d6", x"22d3", x"22d0", 
    x"22cd", x"22ca", x"22c7", x"22c4", x"22c1", x"22be", x"22bb", x"22b8", 
    x"22b5", x"22b2", x"22af", x"22ac", x"22a9", x"22a5", x"22a2", x"229f", 
    x"229c", x"2299", x"2296", x"2293", x"2290", x"228d", x"228a", x"2287", 
    x"2284", x"2281", x"227e", x"227b", x"2278", x"2275", x"2272", x"226f", 
    x"226c", x"2269", x"2266", x"2263", x"2260", x"225d", x"225a", x"2257", 
    x"2254", x"2251", x"224e", x"224b", x"2248", x"2245", x"2242", x"223f", 
    x"223c", x"2239", x"2236", x"2233", x"222f", x"222c", x"2229", x"2226", 
    x"2223", x"2220", x"221d", x"221a", x"2217", x"2214", x"2211", x"220e", 
    x"220b", x"2208", x"2205", x"2202", x"21ff", x"21fc", x"21f9", x"21f6", 
    x"21f3", x"21f0", x"21ed", x"21ea", x"21e7", x"21e4", x"21e1", x"21de", 
    x"21db", x"21d8", x"21d5", x"21d2", x"21cf", x"21cc", x"21c9", x"21c5", 
    x"21c2", x"21bf", x"21bc", x"21b9", x"21b6", x"21b3", x"21b0", x"21ad", 
    x"21aa", x"21a7", x"21a4", x"21a1", x"219e", x"219b", x"2198", x"2195", 
    x"2192", x"218f", x"218c", x"2189", x"2186", x"2183", x"2180", x"217d", 
    x"217a", x"2177", x"2174", x"2171", x"216e", x"216b", x"2168", x"2164", 
    x"2161", x"215e", x"215b", x"2158", x"2155", x"2152", x"214f", x"214c", 
    x"2149", x"2146", x"2143", x"2140", x"213d", x"213a", x"2137", x"2134", 
    x"2131", x"212e", x"212b", x"2128", x"2125", x"2122", x"211f", x"211c", 
    x"2119", x"2116", x"2113", x"2110", x"210c", x"2109", x"2106", x"2103", 
    x"2100", x"20fd", x"20fa", x"20f7", x"20f4", x"20f1", x"20ee", x"20eb", 
    x"20e8", x"20e5", x"20e2", x"20df", x"20dc", x"20d9", x"20d6", x"20d3", 
    x"20d0", x"20cd", x"20ca", x"20c7", x"20c4", x"20c1", x"20be", x"20bb", 
    x"20b7", x"20b4", x"20b1", x"20ae", x"20ab", x"20a8", x"20a5", x"20a2", 
    x"209f", x"209c", x"2099", x"2096", x"2093", x"2090", x"208d", x"208a", 
    x"2087", x"2084", x"2081", x"207e", x"207b", x"2078", x"2075", x"2072", 
    x"206f", x"206c", x"2068", x"2065", x"2062", x"205f", x"205c", x"2059", 
    x"2056", x"2053", x"2050", x"204d", x"204a", x"2047", x"2044", x"2041", 
    x"203e", x"203b", x"2038", x"2035", x"2032", x"202f", x"202c", x"2029", 
    x"2026", x"2023", x"2020", x"201c", x"2019", x"2016", x"2013", x"2010", 
    x"200d", x"200a", x"2007", x"2004", x"2001", x"1ffe", x"1ffb", x"1ff8", 
    x"1ff5", x"1ff2", x"1fef", x"1fec", x"1fe9", x"1fe6", x"1fe3", x"1fe0", 
    x"1fdd", x"1fda", x"1fd7", x"1fd3", x"1fd0", x"1fcd", x"1fca", x"1fc7", 
    x"1fc4", x"1fc1", x"1fbe", x"1fbb", x"1fb8", x"1fb5", x"1fb2", x"1faf", 
    x"1fac", x"1fa9", x"1fa6", x"1fa3", x"1fa0", x"1f9d", x"1f9a", x"1f97", 
    x"1f94", x"1f91", x"1f8d", x"1f8a", x"1f87", x"1f84", x"1f81", x"1f7e", 
    x"1f7b", x"1f78", x"1f75", x"1f72", x"1f6f", x"1f6c", x"1f69", x"1f66", 
    x"1f63", x"1f60", x"1f5d", x"1f5a", x"1f57", x"1f54", x"1f51", x"1f4e", 
    x"1f4a", x"1f47", x"1f44", x"1f41", x"1f3e", x"1f3b", x"1f38", x"1f35", 
    x"1f32", x"1f2f", x"1f2c", x"1f29", x"1f26", x"1f23", x"1f20", x"1f1d", 
    x"1f1a", x"1f17", x"1f14", x"1f11", x"1f0e", x"1f0a", x"1f07", x"1f04", 
    x"1f01", x"1efe", x"1efb", x"1ef8", x"1ef5", x"1ef2", x"1eef", x"1eec", 
    x"1ee9", x"1ee6", x"1ee3", x"1ee0", x"1edd", x"1eda", x"1ed7", x"1ed4", 
    x"1ed1", x"1ece", x"1eca", x"1ec7", x"1ec4", x"1ec1", x"1ebe", x"1ebb", 
    x"1eb8", x"1eb5", x"1eb2", x"1eaf", x"1eac", x"1ea9", x"1ea6", x"1ea3", 
    x"1ea0", x"1e9d", x"1e9a", x"1e97", x"1e94", x"1e91", x"1e8d", x"1e8a", 
    x"1e87", x"1e84", x"1e81", x"1e7e", x"1e7b", x"1e78", x"1e75", x"1e72", 
    x"1e6f", x"1e6c", x"1e69", x"1e66", x"1e63", x"1e60", x"1e5d", x"1e5a", 
    x"1e57", x"1e54", x"1e50", x"1e4d", x"1e4a", x"1e47", x"1e44", x"1e41", 
    x"1e3e", x"1e3b", x"1e38", x"1e35", x"1e32", x"1e2f", x"1e2c", x"1e29", 
    x"1e26", x"1e23", x"1e20", x"1e1d", x"1e19", x"1e16", x"1e13", x"1e10", 
    x"1e0d", x"1e0a", x"1e07", x"1e04", x"1e01", x"1dfe", x"1dfb", x"1df8", 
    x"1df5", x"1df2", x"1def", x"1dec", x"1de9", x"1de6", x"1de3", x"1ddf", 
    x"1ddc", x"1dd9", x"1dd6", x"1dd3", x"1dd0", x"1dcd", x"1dca", x"1dc7", 
    x"1dc4", x"1dc1", x"1dbe", x"1dbb", x"1db8", x"1db5", x"1db2", x"1daf", 
    x"1dac", x"1da8", x"1da5", x"1da2", x"1d9f", x"1d9c", x"1d99", x"1d96", 
    x"1d93", x"1d90", x"1d8d", x"1d8a", x"1d87", x"1d84", x"1d81", x"1d7e", 
    x"1d7b", x"1d78", x"1d75", x"1d71", x"1d6e", x"1d6b", x"1d68", x"1d65", 
    x"1d62", x"1d5f", x"1d5c", x"1d59", x"1d56", x"1d53", x"1d50", x"1d4d", 
    x"1d4a", x"1d47", x"1d44", x"1d41", x"1d3d", x"1d3a", x"1d37", x"1d34", 
    x"1d31", x"1d2e", x"1d2b", x"1d28", x"1d25", x"1d22", x"1d1f", x"1d1c", 
    x"1d19", x"1d16", x"1d13", x"1d10", x"1d0d", x"1d09", x"1d06", x"1d03", 
    x"1d00", x"1cfd", x"1cfa", x"1cf7", x"1cf4", x"1cf1", x"1cee", x"1ceb", 
    x"1ce8", x"1ce5", x"1ce2", x"1cdf", x"1cdc", x"1cd9", x"1cd5", x"1cd2", 
    x"1ccf", x"1ccc", x"1cc9", x"1cc6", x"1cc3", x"1cc0", x"1cbd", x"1cba", 
    x"1cb7", x"1cb4", x"1cb1", x"1cae", x"1cab", x"1ca8", x"1ca4", x"1ca1", 
    x"1c9e", x"1c9b", x"1c98", x"1c95", x"1c92", x"1c8f", x"1c8c", x"1c89", 
    x"1c86", x"1c83", x"1c80", x"1c7d", x"1c7a", x"1c77", x"1c73", x"1c70", 
    x"1c6d", x"1c6a", x"1c67", x"1c64", x"1c61", x"1c5e", x"1c5b", x"1c58", 
    x"1c55", x"1c52", x"1c4f", x"1c4c", x"1c49", x"1c46", x"1c42", x"1c3f", 
    x"1c3c", x"1c39", x"1c36", x"1c33", x"1c30", x"1c2d", x"1c2a", x"1c27", 
    x"1c24", x"1c21", x"1c1e", x"1c1b", x"1c18", x"1c14", x"1c11", x"1c0e", 
    x"1c0b", x"1c08", x"1c05", x"1c02", x"1bff", x"1bfc", x"1bf9", x"1bf6", 
    x"1bf3", x"1bf0", x"1bed", x"1bea", x"1be7", x"1be3", x"1be0", x"1bdd", 
    x"1bda", x"1bd7", x"1bd4", x"1bd1", x"1bce", x"1bcb", x"1bc8", x"1bc5", 
    x"1bc2", x"1bbf", x"1bbc", x"1bb9", x"1bb5", x"1bb2", x"1baf", x"1bac", 
    x"1ba9", x"1ba6", x"1ba3", x"1ba0", x"1b9d", x"1b9a", x"1b97", x"1b94", 
    x"1b91", x"1b8e", x"1b8a", x"1b87", x"1b84", x"1b81", x"1b7e", x"1b7b", 
    x"1b78", x"1b75", x"1b72", x"1b6f", x"1b6c", x"1b69", x"1b66", x"1b63", 
    x"1b60", x"1b5c", x"1b59", x"1b56", x"1b53", x"1b50", x"1b4d", x"1b4a", 
    x"1b47", x"1b44", x"1b41", x"1b3e", x"1b3b", x"1b38", x"1b35", x"1b31", 
    x"1b2e", x"1b2b", x"1b28", x"1b25", x"1b22", x"1b1f", x"1b1c", x"1b19", 
    x"1b16", x"1b13", x"1b10", x"1b0d", x"1b0a", x"1b07", x"1b03", x"1b00", 
    x"1afd", x"1afa", x"1af7", x"1af4", x"1af1", x"1aee", x"1aeb", x"1ae8", 
    x"1ae5", x"1ae2", x"1adf", x"1adc", x"1ad8", x"1ad5", x"1ad2", x"1acf", 
    x"1acc", x"1ac9", x"1ac6", x"1ac3", x"1ac0", x"1abd", x"1aba", x"1ab7", 
    x"1ab4", x"1ab1", x"1aad", x"1aaa", x"1aa7", x"1aa4", x"1aa1", x"1a9e", 
    x"1a9b", x"1a98", x"1a95", x"1a92", x"1a8f", x"1a8c", x"1a89", x"1a85", 
    x"1a82", x"1a7f", x"1a7c", x"1a79", x"1a76", x"1a73", x"1a70", x"1a6d", 
    x"1a6a", x"1a67", x"1a64", x"1a61", x"1a5e", x"1a5a", x"1a57", x"1a54", 
    x"1a51", x"1a4e", x"1a4b", x"1a48", x"1a45", x"1a42", x"1a3f", x"1a3c", 
    x"1a39", x"1a36", x"1a32", x"1a2f", x"1a2c", x"1a29", x"1a26", x"1a23", 
    x"1a20", x"1a1d", x"1a1a", x"1a17", x"1a14", x"1a11", x"1a0e", x"1a0b", 
    x"1a07", x"1a04", x"1a01", x"19fe", x"19fb", x"19f8", x"19f5", x"19f2", 
    x"19ef", x"19ec", x"19e9", x"19e6", x"19e3", x"19df", x"19dc", x"19d9", 
    x"19d6", x"19d3", x"19d0", x"19cd", x"19ca", x"19c7", x"19c4", x"19c1", 
    x"19be", x"19bb", x"19b7", x"19b4", x"19b1", x"19ae", x"19ab", x"19a8", 
    x"19a5", x"19a2", x"199f", x"199c", x"1999", x"1996", x"1993", x"198f", 
    x"198c", x"1989", x"1986", x"1983", x"1980", x"197d", x"197a", x"1977", 
    x"1974", x"1971", x"196e", x"196a", x"1967", x"1964", x"1961", x"195e", 
    x"195b", x"1958", x"1955", x"1952", x"194f", x"194c", x"1949", x"1946", 
    x"1942", x"193f", x"193c", x"1939", x"1936", x"1933", x"1930", x"192d", 
    x"192a", x"1927", x"1924", x"1921", x"191d", x"191a", x"1917", x"1914", 
    x"1911", x"190e", x"190b", x"1908", x"1905", x"1902", x"18ff", x"18fc", 
    x"18f9", x"18f5", x"18f2", x"18ef", x"18ec", x"18e9", x"18e6", x"18e3", 
    x"18e0", x"18dd", x"18da", x"18d7", x"18d4", x"18d0", x"18cd", x"18ca", 
    x"18c7", x"18c4", x"18c1", x"18be", x"18bb", x"18b8", x"18b5", x"18b2", 
    x"18af", x"18ab", x"18a8", x"18a5", x"18a2", x"189f", x"189c", x"1899", 
    x"1896", x"1893", x"1890", x"188d", x"188a", x"1886", x"1883", x"1880", 
    x"187d", x"187a", x"1877", x"1874", x"1871", x"186e", x"186b", x"1868", 
    x"1865", x"1861", x"185e", x"185b", x"1858", x"1855", x"1852", x"184f", 
    x"184c", x"1849", x"1846", x"1843", x"1840", x"183c", x"1839", x"1836", 
    x"1833", x"1830", x"182d", x"182a", x"1827", x"1824", x"1821", x"181e", 
    x"181b", x"1817", x"1814", x"1811", x"180e", x"180b", x"1808", x"1805", 
    x"1802", x"17ff", x"17fc", x"17f9", x"17f6", x"17f2", x"17ef", x"17ec", 
    x"17e9", x"17e6", x"17e3", x"17e0", x"17dd", x"17da", x"17d7", x"17d4", 
    x"17d0", x"17cd", x"17ca", x"17c7", x"17c4", x"17c1", x"17be", x"17bb", 
    x"17b8", x"17b5", x"17b2", x"17af", x"17ab", x"17a8", x"17a5", x"17a2", 
    x"179f", x"179c", x"1799", x"1796", x"1793", x"1790", x"178d", x"1789", 
    x"1786", x"1783", x"1780", x"177d", x"177a", x"1777", x"1774", x"1771", 
    x"176e", x"176b", x"1767", x"1764", x"1761", x"175e", x"175b", x"1758", 
    x"1755", x"1752", x"174f", x"174c", x"1749", x"1746", x"1742", x"173f", 
    x"173c", x"1739", x"1736", x"1733", x"1730", x"172d", x"172a", x"1727", 
    x"1724", x"1720", x"171d", x"171a", x"1717", x"1714", x"1711", x"170e", 
    x"170b", x"1708", x"1705", x"1702", x"16fe", x"16fb", x"16f8", x"16f5", 
    x"16f2", x"16ef", x"16ec", x"16e9", x"16e6", x"16e3", x"16e0", x"16dc", 
    x"16d9", x"16d6", x"16d3", x"16d0", x"16cd", x"16ca", x"16c7", x"16c4", 
    x"16c1", x"16be", x"16ba", x"16b7", x"16b4", x"16b1", x"16ae", x"16ab", 
    x"16a8", x"16a5", x"16a2", x"169f", x"169c", x"1698", x"1695", x"1692", 
    x"168f", x"168c", x"1689", x"1686", x"1683", x"1680", x"167d", x"167a", 
    x"1676", x"1673", x"1670", x"166d", x"166a", x"1667", x"1664", x"1661", 
    x"165e", x"165b", x"1657", x"1654", x"1651", x"164e", x"164b", x"1648", 
    x"1645", x"1642", x"163f", x"163c", x"1639", x"1635", x"1632", x"162f", 
    x"162c", x"1629", x"1626", x"1623", x"1620", x"161d", x"161a", x"1617", 
    x"1613", x"1610", x"160d", x"160a", x"1607", x"1604", x"1601", x"15fe", 
    x"15fb", x"15f8", x"15f4", x"15f1", x"15ee", x"15eb", x"15e8", x"15e5", 
    x"15e2", x"15df", x"15dc", x"15d9", x"15d6", x"15d2", x"15cf", x"15cc", 
    x"15c9", x"15c6", x"15c3", x"15c0", x"15bd", x"15ba", x"15b7", x"15b3", 
    x"15b0", x"15ad", x"15aa", x"15a7", x"15a4", x"15a1", x"159e", x"159b", 
    x"1598", x"1595", x"1591", x"158e", x"158b", x"1588", x"1585", x"1582", 
    x"157f", x"157c", x"1579", x"1576", x"1572", x"156f", x"156c", x"1569", 
    x"1566", x"1563", x"1560", x"155d", x"155a", x"1557", x"1553", x"1550", 
    x"154d", x"154a", x"1547", x"1544", x"1541", x"153e", x"153b", x"1538", 
    x"1534", x"1531", x"152e", x"152b", x"1528", x"1525", x"1522", x"151f", 
    x"151c", x"1519", x"1516", x"1512", x"150f", x"150c", x"1509", x"1506", 
    x"1503", x"1500", x"14fd", x"14fa", x"14f7", x"14f3", x"14f0", x"14ed", 
    x"14ea", x"14e7", x"14e4", x"14e1", x"14de", x"14db", x"14d8", x"14d4", 
    x"14d1", x"14ce", x"14cb", x"14c8", x"14c5", x"14c2", x"14bf", x"14bc", 
    x"14b9", x"14b5", x"14b2", x"14af", x"14ac", x"14a9", x"14a6", x"14a3", 
    x"14a0", x"149d", x"149a", x"1496", x"1493", x"1490", x"148d", x"148a", 
    x"1487", x"1484", x"1481", x"147e", x"147b", x"1477", x"1474", x"1471", 
    x"146e", x"146b", x"1468", x"1465", x"1462", x"145f", x"145c", x"1458", 
    x"1455", x"1452", x"144f", x"144c", x"1449", x"1446", x"1443", x"1440", 
    x"143c", x"1439", x"1436", x"1433", x"1430", x"142d", x"142a", x"1427", 
    x"1424", x"1421", x"141d", x"141a", x"1417", x"1414", x"1411", x"140e", 
    x"140b", x"1408", x"1405", x"1402", x"13fe", x"13fb", x"13f8", x"13f5", 
    x"13f2", x"13ef", x"13ec", x"13e9", x"13e6", x"13e3", x"13df", x"13dc", 
    x"13d9", x"13d6", x"13d3", x"13d0", x"13cd", x"13ca", x"13c7", x"13c3", 
    x"13c0", x"13bd", x"13ba", x"13b7", x"13b4", x"13b1", x"13ae", x"13ab", 
    x"13a8", x"13a4", x"13a1", x"139e", x"139b", x"1398", x"1395", x"1392", 
    x"138f", x"138c", x"1388", x"1385", x"1382", x"137f", x"137c", x"1379", 
    x"1376", x"1373", x"1370", x"136d", x"1369", x"1366", x"1363", x"1360", 
    x"135d", x"135a", x"1357", x"1354", x"1351", x"134d", x"134a", x"1347", 
    x"1344", x"1341", x"133e", x"133b", x"1338", x"1335", x"1332", x"132e", 
    x"132b", x"1328", x"1325", x"1322", x"131f", x"131c", x"1319", x"1316", 
    x"1312", x"130f", x"130c", x"1309", x"1306", x"1303", x"1300", x"12fd", 
    x"12fa", x"12f7", x"12f3", x"12f0", x"12ed", x"12ea", x"12e7", x"12e4", 
    x"12e1", x"12de", x"12db", x"12d7", x"12d4", x"12d1", x"12ce", x"12cb", 
    x"12c8", x"12c5", x"12c2", x"12bf", x"12bb", x"12b8", x"12b5", x"12b2", 
    x"12af", x"12ac", x"12a9", x"12a6", x"12a3", x"12a0", x"129c", x"1299", 
    x"1296", x"1293", x"1290", x"128d", x"128a", x"1287", x"1284", x"1280", 
    x"127d", x"127a", x"1277", x"1274", x"1271", x"126e", x"126b", x"1268", 
    x"1264", x"1261", x"125e", x"125b", x"1258", x"1255", x"1252", x"124f", 
    x"124c", x"1248", x"1245", x"1242", x"123f", x"123c", x"1239", x"1236", 
    x"1233", x"1230", x"122c", x"1229", x"1226", x"1223", x"1220", x"121d", 
    x"121a", x"1217", x"1214", x"1210", x"120d", x"120a", x"1207", x"1204", 
    x"1201", x"11fe", x"11fb", x"11f8", x"11f5", x"11f1", x"11ee", x"11eb", 
    x"11e8", x"11e5", x"11e2", x"11df", x"11dc", x"11d9", x"11d5", x"11d2", 
    x"11cf", x"11cc", x"11c9", x"11c6", x"11c3", x"11c0", x"11bd", x"11b9", 
    x"11b6", x"11b3", x"11b0", x"11ad", x"11aa", x"11a7", x"11a4", x"11a1", 
    x"119d", x"119a", x"1197", x"1194", x"1191", x"118e", x"118b", x"1188", 
    x"1185", x"1181", x"117e", x"117b", x"1178", x"1175", x"1172", x"116f", 
    x"116c", x"1168", x"1165", x"1162", x"115f", x"115c", x"1159", x"1156", 
    x"1153", x"1150", x"114c", x"1149", x"1146", x"1143", x"1140", x"113d", 
    x"113a", x"1137", x"1134", x"1130", x"112d", x"112a", x"1127", x"1124", 
    x"1121", x"111e", x"111b", x"1118", x"1114", x"1111", x"110e", x"110b", 
    x"1108", x"1105", x"1102", x"10ff", x"10fc", x"10f8", x"10f5", x"10f2", 
    x"10ef", x"10ec", x"10e9", x"10e6", x"10e3", x"10e0", x"10dc", x"10d9", 
    x"10d6", x"10d3", x"10d0", x"10cd", x"10ca", x"10c7", x"10c3", x"10c0", 
    x"10bd", x"10ba", x"10b7", x"10b4", x"10b1", x"10ae", x"10ab", x"10a7", 
    x"10a4", x"10a1", x"109e", x"109b", x"1098", x"1095", x"1092", x"108f", 
    x"108b", x"1088", x"1085", x"1082", x"107f", x"107c", x"1079", x"1076", 
    x"1072", x"106f", x"106c", x"1069", x"1066", x"1063", x"1060", x"105d", 
    x"105a", x"1056", x"1053", x"1050", x"104d", x"104a", x"1047", x"1044", 
    x"1041", x"103e", x"103a", x"1037", x"1034", x"1031", x"102e", x"102b", 
    x"1028", x"1025", x"1021", x"101e", x"101b", x"1018", x"1015", x"1012", 
    x"100f", x"100c", x"1009", x"1005", x"1002", x"0fff", x"0ffc", x"0ff9", 
    x"0ff6", x"0ff3", x"0ff0", x"0fec", x"0fe9", x"0fe6", x"0fe3", x"0fe0", 
    x"0fdd", x"0fda", x"0fd7", x"0fd4", x"0fd0", x"0fcd", x"0fca", x"0fc7", 
    x"0fc4", x"0fc1", x"0fbe", x"0fbb", x"0fb8", x"0fb4", x"0fb1", x"0fae", 
    x"0fab", x"0fa8", x"0fa5", x"0fa2", x"0f9f", x"0f9b", x"0f98", x"0f95", 
    x"0f92", x"0f8f", x"0f8c", x"0f89", x"0f86", x"0f82", x"0f7f", x"0f7c", 
    x"0f79", x"0f76", x"0f73", x"0f70", x"0f6d", x"0f6a", x"0f66", x"0f63", 
    x"0f60", x"0f5d", x"0f5a", x"0f57", x"0f54", x"0f51", x"0f4d", x"0f4a", 
    x"0f47", x"0f44", x"0f41", x"0f3e", x"0f3b", x"0f38", x"0f35", x"0f31", 
    x"0f2e", x"0f2b", x"0f28", x"0f25", x"0f22", x"0f1f", x"0f1c", x"0f18", 
    x"0f15", x"0f12", x"0f0f", x"0f0c", x"0f09", x"0f06", x"0f03", x"0eff", 
    x"0efc", x"0ef9", x"0ef6", x"0ef3", x"0ef0", x"0eed", x"0eea", x"0ee7", 
    x"0ee3", x"0ee0", x"0edd", x"0eda", x"0ed7", x"0ed4", x"0ed1", x"0ece", 
    x"0eca", x"0ec7", x"0ec4", x"0ec1", x"0ebe", x"0ebb", x"0eb8", x"0eb5", 
    x"0eb1", x"0eae", x"0eab", x"0ea8", x"0ea5", x"0ea2", x"0e9f", x"0e9c", 
    x"0e99", x"0e95", x"0e92", x"0e8f", x"0e8c", x"0e89", x"0e86", x"0e83", 
    x"0e80", x"0e7c", x"0e79", x"0e76", x"0e73", x"0e70", x"0e6d", x"0e6a", 
    x"0e67", x"0e63", x"0e60", x"0e5d", x"0e5a", x"0e57", x"0e54", x"0e51", 
    x"0e4e", x"0e4a", x"0e47", x"0e44", x"0e41", x"0e3e", x"0e3b", x"0e38", 
    x"0e35", x"0e32", x"0e2e", x"0e2b", x"0e28", x"0e25", x"0e22", x"0e1f", 
    x"0e1c", x"0e19", x"0e15", x"0e12", x"0e0f", x"0e0c", x"0e09", x"0e06", 
    x"0e03", x"0e00", x"0dfc", x"0df9", x"0df6", x"0df3", x"0df0", x"0ded", 
    x"0dea", x"0de7", x"0de3", x"0de0", x"0ddd", x"0dda", x"0dd7", x"0dd4", 
    x"0dd1", x"0dce", x"0dca", x"0dc7", x"0dc4", x"0dc1", x"0dbe", x"0dbb", 
    x"0db8", x"0db5", x"0db1", x"0dae", x"0dab", x"0da8", x"0da5", x"0da2", 
    x"0d9f", x"0d9c", x"0d98", x"0d95", x"0d92", x"0d8f", x"0d8c", x"0d89", 
    x"0d86", x"0d83", x"0d7f", x"0d7c", x"0d79", x"0d76", x"0d73", x"0d70", 
    x"0d6d", x"0d6a", x"0d66", x"0d63", x"0d60", x"0d5d", x"0d5a", x"0d57", 
    x"0d54", x"0d51", x"0d4e", x"0d4a", x"0d47", x"0d44", x"0d41", x"0d3e", 
    x"0d3b", x"0d38", x"0d35", x"0d31", x"0d2e", x"0d2b", x"0d28", x"0d25", 
    x"0d22", x"0d1f", x"0d1c", x"0d18", x"0d15", x"0d12", x"0d0f", x"0d0c", 
    x"0d09", x"0d06", x"0d03", x"0cff", x"0cfc", x"0cf9", x"0cf6", x"0cf3", 
    x"0cf0", x"0ced", x"0cea", x"0ce6", x"0ce3", x"0ce0", x"0cdd", x"0cda", 
    x"0cd7", x"0cd4", x"0cd1", x"0ccd", x"0cca", x"0cc7", x"0cc4", x"0cc1", 
    x"0cbe", x"0cbb", x"0cb7", x"0cb4", x"0cb1", x"0cae", x"0cab", x"0ca8", 
    x"0ca5", x"0ca2", x"0c9e", x"0c9b", x"0c98", x"0c95", x"0c92", x"0c8f", 
    x"0c8c", x"0c89", x"0c85", x"0c82", x"0c7f", x"0c7c", x"0c79", x"0c76", 
    x"0c73", x"0c70", x"0c6c", x"0c69", x"0c66", x"0c63", x"0c60", x"0c5d", 
    x"0c5a", x"0c57", x"0c53", x"0c50", x"0c4d", x"0c4a", x"0c47", x"0c44", 
    x"0c41", x"0c3e", x"0c3a", x"0c37", x"0c34", x"0c31", x"0c2e", x"0c2b", 
    x"0c28", x"0c25", x"0c21", x"0c1e", x"0c1b", x"0c18", x"0c15", x"0c12", 
    x"0c0f", x"0c0c", x"0c08", x"0c05", x"0c02", x"0bff", x"0bfc", x"0bf9", 
    x"0bf6", x"0bf3", x"0bef", x"0bec", x"0be9", x"0be6", x"0be3", x"0be0", 
    x"0bdd", x"0bd9", x"0bd6", x"0bd3", x"0bd0", x"0bcd", x"0bca", x"0bc7", 
    x"0bc4", x"0bc0", x"0bbd", x"0bba", x"0bb7", x"0bb4", x"0bb1", x"0bae", 
    x"0bab", x"0ba7", x"0ba4", x"0ba1", x"0b9e", x"0b9b", x"0b98", x"0b95", 
    x"0b92", x"0b8e", x"0b8b", x"0b88", x"0b85", x"0b82", x"0b7f", x"0b7c", 
    x"0b78", x"0b75", x"0b72", x"0b6f", x"0b6c", x"0b69", x"0b66", x"0b63", 
    x"0b5f", x"0b5c", x"0b59", x"0b56", x"0b53", x"0b50", x"0b4d", x"0b4a", 
    x"0b46", x"0b43", x"0b40", x"0b3d", x"0b3a", x"0b37", x"0b34", x"0b31", 
    x"0b2d", x"0b2a", x"0b27", x"0b24", x"0b21", x"0b1e", x"0b1b", x"0b17", 
    x"0b14", x"0b11", x"0b0e", x"0b0b", x"0b08", x"0b05", x"0b02", x"0afe", 
    x"0afb", x"0af8", x"0af5", x"0af2", x"0aef", x"0aec", x"0ae9", x"0ae5", 
    x"0ae2", x"0adf", x"0adc", x"0ad9", x"0ad6", x"0ad3", x"0acf", x"0acc", 
    x"0ac9", x"0ac6", x"0ac3", x"0ac0", x"0abd", x"0aba", x"0ab6", x"0ab3", 
    x"0ab0", x"0aad", x"0aaa", x"0aa7", x"0aa4", x"0aa1", x"0a9d", x"0a9a", 
    x"0a97", x"0a94", x"0a91", x"0a8e", x"0a8b", x"0a87", x"0a84", x"0a81", 
    x"0a7e", x"0a7b", x"0a78", x"0a75", x"0a72", x"0a6e", x"0a6b", x"0a68", 
    x"0a65", x"0a62", x"0a5f", x"0a5c", x"0a59", x"0a55", x"0a52", x"0a4f", 
    x"0a4c", x"0a49", x"0a46", x"0a43", x"0a3f", x"0a3c", x"0a39", x"0a36", 
    x"0a33", x"0a30", x"0a2d", x"0a2a", x"0a26", x"0a23", x"0a20", x"0a1d", 
    x"0a1a", x"0a17", x"0a14", x"0a11", x"0a0d", x"0a0a", x"0a07", x"0a04", 
    x"0a01", x"09fe", x"09fb", x"09f7", x"09f4", x"09f1", x"09ee", x"09eb", 
    x"09e8", x"09e5", x"09e2", x"09de", x"09db", x"09d8", x"09d5", x"09d2", 
    x"09cf", x"09cc", x"09c8", x"09c5", x"09c2", x"09bf", x"09bc", x"09b9", 
    x"09b6", x"09b3", x"09af", x"09ac", x"09a9", x"09a6", x"09a3", x"09a0", 
    x"099d", x"0999", x"0996", x"0993", x"0990", x"098d", x"098a", x"0987", 
    x"0984", x"0980", x"097d", x"097a", x"0977", x"0974", x"0971", x"096e", 
    x"096a", x"0967", x"0964", x"0961", x"095e", x"095b", x"0958", x"0955", 
    x"0951", x"094e", x"094b", x"0948", x"0945", x"0942", x"093f", x"093b", 
    x"0938", x"0935", x"0932", x"092f", x"092c", x"0929", x"0926", x"0922", 
    x"091f", x"091c", x"0919", x"0916", x"0913", x"0910", x"090c", x"0909", 
    x"0906", x"0903", x"0900", x"08fd", x"08fa", x"08f7", x"08f3", x"08f0", 
    x"08ed", x"08ea", x"08e7", x"08e4", x"08e1", x"08dd", x"08da", x"08d7", 
    x"08d4", x"08d1", x"08ce", x"08cb", x"08c8", x"08c4", x"08c1", x"08be", 
    x"08bb", x"08b8", x"08b5", x"08b2", x"08ae", x"08ab", x"08a8", x"08a5", 
    x"08a2", x"089f", x"089c", x"0899", x"0895", x"0892", x"088f", x"088c", 
    x"0889", x"0886", x"0883", x"087f", x"087c", x"0879", x"0876", x"0873", 
    x"0870", x"086d", x"086a", x"0866", x"0863", x"0860", x"085d", x"085a", 
    x"0857", x"0854", x"0850", x"084d", x"084a", x"0847", x"0844", x"0841", 
    x"083e", x"083a", x"0837", x"0834", x"0831", x"082e", x"082b", x"0828", 
    x"0825", x"0821", x"081e", x"081b", x"0818", x"0815", x"0812", x"080f", 
    x"080b", x"0808", x"0805", x"0802", x"07ff", x"07fc", x"07f9", x"07f6", 
    x"07f2", x"07ef", x"07ec", x"07e9", x"07e6", x"07e3", x"07e0", x"07dc", 
    x"07d9", x"07d6", x"07d3", x"07d0", x"07cd", x"07ca", x"07c6", x"07c3", 
    x"07c0", x"07bd", x"07ba", x"07b7", x"07b4", x"07b1", x"07ad", x"07aa", 
    x"07a7", x"07a4", x"07a1", x"079e", x"079b", x"0797", x"0794", x"0791", 
    x"078e", x"078b", x"0788", x"0785", x"0781", x"077e", x"077b", x"0778", 
    x"0775", x"0772", x"076f", x"076c", x"0768", x"0765", x"0762", x"075f", 
    x"075c", x"0759", x"0756", x"0752", x"074f", x"074c", x"0749", x"0746", 
    x"0743", x"0740", x"073c", x"0739", x"0736", x"0733", x"0730", x"072d", 
    x"072a", x"0727", x"0723", x"0720", x"071d", x"071a", x"0717", x"0714", 
    x"0711", x"070d", x"070a", x"0707", x"0704", x"0701", x"06fe", x"06fb", 
    x"06f7", x"06f4", x"06f1", x"06ee", x"06eb", x"06e8", x"06e5", x"06e2", 
    x"06de", x"06db", x"06d8", x"06d5", x"06d2", x"06cf", x"06cc", x"06c8", 
    x"06c5", x"06c2", x"06bf", x"06bc", x"06b9", x"06b6", x"06b2", x"06af", 
    x"06ac", x"06a9", x"06a6", x"06a3", x"06a0", x"069d", x"0699", x"0696", 
    x"0693", x"0690", x"068d", x"068a", x"0687", x"0683", x"0680", x"067d", 
    x"067a", x"0677", x"0674", x"0671", x"066d", x"066a", x"0667", x"0664", 
    x"0661", x"065e", x"065b", x"0657", x"0654", x"0651", x"064e", x"064b", 
    x"0648", x"0645", x"0642", x"063e", x"063b", x"0638", x"0635", x"0632", 
    x"062f", x"062c", x"0628", x"0625", x"0622", x"061f", x"061c", x"0619", 
    x"0616", x"0612", x"060f", x"060c", x"0609", x"0606", x"0603", x"0600", 
    x"05fc", x"05f9", x"05f6", x"05f3", x"05f0", x"05ed", x"05ea", x"05e7", 
    x"05e3", x"05e0", x"05dd", x"05da", x"05d7", x"05d4", x"05d1", x"05cd", 
    x"05ca", x"05c7", x"05c4", x"05c1", x"05be", x"05bb", x"05b7", x"05b4", 
    x"05b1", x"05ae", x"05ab", x"05a8", x"05a5", x"05a1", x"059e", x"059b", 
    x"0598", x"0595", x"0592", x"058f", x"058c", x"0588", x"0585", x"0582", 
    x"057f", x"057c", x"0579", x"0576", x"0572", x"056f", x"056c", x"0569", 
    x"0566", x"0563", x"0560", x"055c", x"0559", x"0556", x"0553", x"0550", 
    x"054d", x"054a", x"0546", x"0543", x"0540", x"053d", x"053a", x"0537", 
    x"0534", x"0530", x"052d", x"052a", x"0527", x"0524", x"0521", x"051e", 
    x"051b", x"0517", x"0514", x"0511", x"050e", x"050b", x"0508", x"0505", 
    x"0501", x"04fe", x"04fb", x"04f8", x"04f5", x"04f2", x"04ef", x"04eb", 
    x"04e8", x"04e5", x"04e2", x"04df", x"04dc", x"04d9", x"04d5", x"04d2", 
    x"04cf", x"04cc", x"04c9", x"04c6", x"04c3", x"04bf", x"04bc", x"04b9", 
    x"04b6", x"04b3", x"04b0", x"04ad", x"04aa", x"04a6", x"04a3", x"04a0", 
    x"049d", x"049a", x"0497", x"0494", x"0490", x"048d", x"048a", x"0487", 
    x"0484", x"0481", x"047e", x"047a", x"0477", x"0474", x"0471", x"046e", 
    x"046b", x"0468", x"0464", x"0461", x"045e", x"045b", x"0458", x"0455", 
    x"0452", x"044e", x"044b", x"0448", x"0445", x"0442", x"043f", x"043c", 
    x"0438", x"0435", x"0432", x"042f", x"042c", x"0429", x"0426", x"0423", 
    x"041f", x"041c", x"0419", x"0416", x"0413", x"0410", x"040d", x"0409", 
    x"0406", x"0403", x"0400", x"03fd", x"03fa", x"03f7", x"03f3", x"03f0", 
    x"03ed", x"03ea", x"03e7", x"03e4", x"03e1", x"03dd", x"03da", x"03d7", 
    x"03d4", x"03d1", x"03ce", x"03cb", x"03c7", x"03c4", x"03c1", x"03be", 
    x"03bb", x"03b8", x"03b5", x"03b1", x"03ae", x"03ab", x"03a8", x"03a5", 
    x"03a2", x"039f", x"039b", x"0398", x"0395", x"0392", x"038f", x"038c", 
    x"0389", x"0385", x"0382", x"037f", x"037c", x"0379", x"0376", x"0373", 
    x"0370", x"036c", x"0369", x"0366", x"0363", x"0360", x"035d", x"035a", 
    x"0356", x"0353", x"0350", x"034d", x"034a", x"0347", x"0344", x"0340", 
    x"033d", x"033a", x"0337", x"0334", x"0331", x"032e", x"032a", x"0327", 
    x"0324", x"0321", x"031e", x"031b", x"0318", x"0314", x"0311", x"030e", 
    x"030b", x"0308", x"0305", x"0302", x"02fe", x"02fb", x"02f8", x"02f5", 
    x"02f2", x"02ef", x"02ec", x"02e8", x"02e5", x"02e2", x"02df", x"02dc", 
    x"02d9", x"02d6", x"02d2", x"02cf", x"02cc", x"02c9", x"02c6", x"02c3", 
    x"02c0", x"02bd", x"02b9", x"02b6", x"02b3", x"02b0", x"02ad", x"02aa", 
    x"02a7", x"02a3", x"02a0", x"029d", x"029a", x"0297", x"0294", x"0291", 
    x"028d", x"028a", x"0287", x"0284", x"0281", x"027e", x"027b", x"0277", 
    x"0274", x"0271", x"026e", x"026b", x"0268", x"0265", x"0261", x"025e", 
    x"025b", x"0258", x"0255", x"0252", x"024f", x"024b", x"0248", x"0245", 
    x"0242", x"023f", x"023c", x"0239", x"0235", x"0232", x"022f", x"022c", 
    x"0229", x"0226", x"0223", x"021f", x"021c", x"0219", x"0216", x"0213", 
    x"0210", x"020d", x"0209", x"0206", x"0203", x"0200", x"01fd", x"01fa", 
    x"01f7", x"01f3", x"01f0", x"01ed", x"01ea", x"01e7", x"01e4", x"01e1", 
    x"01dd", x"01da", x"01d7", x"01d4", x"01d1", x"01ce", x"01cb", x"01c8", 
    x"01c4", x"01c1", x"01be", x"01bb", x"01b8", x"01b5", x"01b2", x"01ae", 
    x"01ab", x"01a8", x"01a5", x"01a2", x"019f", x"019c", x"0198", x"0195", 
    x"0192", x"018f", x"018c", x"0189", x"0186", x"0182", x"017f", x"017c", 
    x"0179", x"0176", x"0173", x"0170", x"016c", x"0169", x"0166", x"0163", 
    x"0160", x"015d", x"015a", x"0156", x"0153", x"0150", x"014d", x"014a", 
    x"0147", x"0144", x"0140", x"013d", x"013a", x"0137", x"0134", x"0131", 
    x"012e", x"012a", x"0127", x"0124", x"0121", x"011e", x"011b", x"0118", 
    x"0114", x"0111", x"010e", x"010b", x"0108", x"0105", x"0102", x"00fe", 
    x"00fb", x"00f8", x"00f5", x"00f2", x"00ef", x"00ec", x"00e8", x"00e5", 
    x"00e2", x"00df", x"00dc", x"00d9", x"00d6", x"00d2", x"00cf", x"00cc", 
    x"00c9", x"00c6", x"00c3", x"00c0", x"00bc", x"00b9", x"00b6", x"00b3", 
    x"00b0", x"00ad", x"00aa", x"00a6", x"00a3", x"00a0", x"009d", x"009a", 
    x"0097", x"0094", x"0091", x"008d", x"008a", x"0087", x"0084", x"0081", 
    x"007e", x"007b", x"0077", x"0074", x"0071", x"006e", x"006b", x"0068", 
    x"0065", x"0061", x"005e", x"005b", x"0058", x"0055", x"0052", x"004f", 
    x"004b", x"0048", x"0045", x"0042", x"003f", x"003c", x"0039", x"0035", 
    x"0032", x"002f", x"002c", x"0029", x"0026", x"0023", x"001f", x"001c", 
    x"0019", x"0016", x"0013", x"0010", x"000d", x"0009", x"0006", x"0003", 
    x"0000", x"fffd", x"fffa", x"fff7", x"fff3", x"fff0", x"ffed", x"ffea", 
    x"ffe7", x"ffe4", x"ffe1", x"ffdd", x"ffda", x"ffd7", x"ffd4", x"ffd1", 
    x"ffce", x"ffcb", x"ffc7", x"ffc4", x"ffc1", x"ffbe", x"ffbb", x"ffb8", 
    x"ffb5", x"ffb1", x"ffae", x"ffab", x"ffa8", x"ffa5", x"ffa2", x"ff9f", 
    x"ff9b", x"ff98", x"ff95", x"ff92", x"ff8f", x"ff8c", x"ff89", x"ff85", 
    x"ff82", x"ff7f", x"ff7c", x"ff79", x"ff76", x"ff73", x"ff6f", x"ff6c", 
    x"ff69", x"ff66", x"ff63", x"ff60", x"ff5d", x"ff5a", x"ff56", x"ff53", 
    x"ff50", x"ff4d", x"ff4a", x"ff47", x"ff44", x"ff40", x"ff3d", x"ff3a", 
    x"ff37", x"ff34", x"ff31", x"ff2e", x"ff2a", x"ff27", x"ff24", x"ff21", 
    x"ff1e", x"ff1b", x"ff18", x"ff14", x"ff11", x"ff0e", x"ff0b", x"ff08", 
    x"ff05", x"ff02", x"fefe", x"fefb", x"fef8", x"fef5", x"fef2", x"feef", 
    x"feec", x"fee8", x"fee5", x"fee2", x"fedf", x"fedc", x"fed9", x"fed6", 
    x"fed2", x"fecf", x"fecc", x"fec9", x"fec6", x"fec3", x"fec0", x"febc", 
    x"feb9", x"feb6", x"feb3", x"feb0", x"fead", x"feaa", x"fea6", x"fea3", 
    x"fea0", x"fe9d", x"fe9a", x"fe97", x"fe94", x"fe90", x"fe8d", x"fe8a", 
    x"fe87", x"fe84", x"fe81", x"fe7e", x"fe7a", x"fe77", x"fe74", x"fe71", 
    x"fe6e", x"fe6b", x"fe68", x"fe64", x"fe61", x"fe5e", x"fe5b", x"fe58", 
    x"fe55", x"fe52", x"fe4e", x"fe4b", x"fe48", x"fe45", x"fe42", x"fe3f", 
    x"fe3c", x"fe38", x"fe35", x"fe32", x"fe2f", x"fe2c", x"fe29", x"fe26", 
    x"fe23", x"fe1f", x"fe1c", x"fe19", x"fe16", x"fe13", x"fe10", x"fe0d", 
    x"fe09", x"fe06", x"fe03", x"fe00", x"fdfd", x"fdfa", x"fdf7", x"fdf3", 
    x"fdf0", x"fded", x"fdea", x"fde7", x"fde4", x"fde1", x"fddd", x"fdda", 
    x"fdd7", x"fdd4", x"fdd1", x"fdce", x"fdcb", x"fdc7", x"fdc4", x"fdc1", 
    x"fdbe", x"fdbb", x"fdb8", x"fdb5", x"fdb1", x"fdae", x"fdab", x"fda8", 
    x"fda5", x"fda2", x"fd9f", x"fd9b", x"fd98", x"fd95", x"fd92", x"fd8f", 
    x"fd8c", x"fd89", x"fd85", x"fd82", x"fd7f", x"fd7c", x"fd79", x"fd76", 
    x"fd73", x"fd6f", x"fd6c", x"fd69", x"fd66", x"fd63", x"fd60", x"fd5d", 
    x"fd59", x"fd56", x"fd53", x"fd50", x"fd4d", x"fd4a", x"fd47", x"fd43", 
    x"fd40", x"fd3d", x"fd3a", x"fd37", x"fd34", x"fd31", x"fd2e", x"fd2a", 
    x"fd27", x"fd24", x"fd21", x"fd1e", x"fd1b", x"fd18", x"fd14", x"fd11", 
    x"fd0e", x"fd0b", x"fd08", x"fd05", x"fd02", x"fcfe", x"fcfb", x"fcf8", 
    x"fcf5", x"fcf2", x"fcef", x"fcec", x"fce8", x"fce5", x"fce2", x"fcdf", 
    x"fcdc", x"fcd9", x"fcd6", x"fcd2", x"fccf", x"fccc", x"fcc9", x"fcc6", 
    x"fcc3", x"fcc0", x"fcbc", x"fcb9", x"fcb6", x"fcb3", x"fcb0", x"fcad", 
    x"fcaa", x"fca6", x"fca3", x"fca0", x"fc9d", x"fc9a", x"fc97", x"fc94", 
    x"fc90", x"fc8d", x"fc8a", x"fc87", x"fc84", x"fc81", x"fc7e", x"fc7b", 
    x"fc77", x"fc74", x"fc71", x"fc6e", x"fc6b", x"fc68", x"fc65", x"fc61", 
    x"fc5e", x"fc5b", x"fc58", x"fc55", x"fc52", x"fc4f", x"fc4b", x"fc48", 
    x"fc45", x"fc42", x"fc3f", x"fc3c", x"fc39", x"fc35", x"fc32", x"fc2f", 
    x"fc2c", x"fc29", x"fc26", x"fc23", x"fc1f", x"fc1c", x"fc19", x"fc16", 
    x"fc13", x"fc10", x"fc0d", x"fc09", x"fc06", x"fc03", x"fc00", x"fbfd", 
    x"fbfa", x"fbf7", x"fbf3", x"fbf0", x"fbed", x"fbea", x"fbe7", x"fbe4", 
    x"fbe1", x"fbdd", x"fbda", x"fbd7", x"fbd4", x"fbd1", x"fbce", x"fbcb", 
    x"fbc8", x"fbc4", x"fbc1", x"fbbe", x"fbbb", x"fbb8", x"fbb5", x"fbb2", 
    x"fbae", x"fbab", x"fba8", x"fba5", x"fba2", x"fb9f", x"fb9c", x"fb98", 
    x"fb95", x"fb92", x"fb8f", x"fb8c", x"fb89", x"fb86", x"fb82", x"fb7f", 
    x"fb7c", x"fb79", x"fb76", x"fb73", x"fb70", x"fb6c", x"fb69", x"fb66", 
    x"fb63", x"fb60", x"fb5d", x"fb5a", x"fb56", x"fb53", x"fb50", x"fb4d", 
    x"fb4a", x"fb47", x"fb44", x"fb41", x"fb3d", x"fb3a", x"fb37", x"fb34", 
    x"fb31", x"fb2e", x"fb2b", x"fb27", x"fb24", x"fb21", x"fb1e", x"fb1b", 
    x"fb18", x"fb15", x"fb11", x"fb0e", x"fb0b", x"fb08", x"fb05", x"fb02", 
    x"faff", x"fafb", x"faf8", x"faf5", x"faf2", x"faef", x"faec", x"fae9", 
    x"fae5", x"fae2", x"fadf", x"fadc", x"fad9", x"fad6", x"fad3", x"fad0", 
    x"facc", x"fac9", x"fac6", x"fac3", x"fac0", x"fabd", x"faba", x"fab6", 
    x"fab3", x"fab0", x"faad", x"faaa", x"faa7", x"faa4", x"faa0", x"fa9d", 
    x"fa9a", x"fa97", x"fa94", x"fa91", x"fa8e", x"fa8a", x"fa87", x"fa84", 
    x"fa81", x"fa7e", x"fa7b", x"fa78", x"fa74", x"fa71", x"fa6e", x"fa6b", 
    x"fa68", x"fa65", x"fa62", x"fa5f", x"fa5b", x"fa58", x"fa55", x"fa52", 
    x"fa4f", x"fa4c", x"fa49", x"fa45", x"fa42", x"fa3f", x"fa3c", x"fa39", 
    x"fa36", x"fa33", x"fa2f", x"fa2c", x"fa29", x"fa26", x"fa23", x"fa20", 
    x"fa1d", x"fa19", x"fa16", x"fa13", x"fa10", x"fa0d", x"fa0a", x"fa07", 
    x"fa04", x"fa00", x"f9fd", x"f9fa", x"f9f7", x"f9f4", x"f9f1", x"f9ee", 
    x"f9ea", x"f9e7", x"f9e4", x"f9e1", x"f9de", x"f9db", x"f9d8", x"f9d4", 
    x"f9d1", x"f9ce", x"f9cb", x"f9c8", x"f9c5", x"f9c2", x"f9be", x"f9bb", 
    x"f9b8", x"f9b5", x"f9b2", x"f9af", x"f9ac", x"f9a9", x"f9a5", x"f9a2", 
    x"f99f", x"f99c", x"f999", x"f996", x"f993", x"f98f", x"f98c", x"f989", 
    x"f986", x"f983", x"f980", x"f97d", x"f979", x"f976", x"f973", x"f970", 
    x"f96d", x"f96a", x"f967", x"f963", x"f960", x"f95d", x"f95a", x"f957", 
    x"f954", x"f951", x"f94e", x"f94a", x"f947", x"f944", x"f941", x"f93e", 
    x"f93b", x"f938", x"f934", x"f931", x"f92e", x"f92b", x"f928", x"f925", 
    x"f922", x"f91e", x"f91b", x"f918", x"f915", x"f912", x"f90f", x"f90c", 
    x"f909", x"f905", x"f902", x"f8ff", x"f8fc", x"f8f9", x"f8f6", x"f8f3", 
    x"f8ef", x"f8ec", x"f8e9", x"f8e6", x"f8e3", x"f8e0", x"f8dd", x"f8d9", 
    x"f8d6", x"f8d3", x"f8d0", x"f8cd", x"f8ca", x"f8c7", x"f8c4", x"f8c0", 
    x"f8bd", x"f8ba", x"f8b7", x"f8b4", x"f8b1", x"f8ae", x"f8aa", x"f8a7", 
    x"f8a4", x"f8a1", x"f89e", x"f89b", x"f898", x"f894", x"f891", x"f88e", 
    x"f88b", x"f888", x"f885", x"f882", x"f87f", x"f87b", x"f878", x"f875", 
    x"f872", x"f86f", x"f86c", x"f869", x"f865", x"f862", x"f85f", x"f85c", 
    x"f859", x"f856", x"f853", x"f84f", x"f84c", x"f849", x"f846", x"f843", 
    x"f840", x"f83d", x"f83a", x"f836", x"f833", x"f830", x"f82d", x"f82a", 
    x"f827", x"f824", x"f820", x"f81d", x"f81a", x"f817", x"f814", x"f811", 
    x"f80e", x"f80a", x"f807", x"f804", x"f801", x"f7fe", x"f7fb", x"f7f8", 
    x"f7f5", x"f7f1", x"f7ee", x"f7eb", x"f7e8", x"f7e5", x"f7e2", x"f7df", 
    x"f7db", x"f7d8", x"f7d5", x"f7d2", x"f7cf", x"f7cc", x"f7c9", x"f7c6", 
    x"f7c2", x"f7bf", x"f7bc", x"f7b9", x"f7b6", x"f7b3", x"f7b0", x"f7ac", 
    x"f7a9", x"f7a6", x"f7a3", x"f7a0", x"f79d", x"f79a", x"f796", x"f793", 
    x"f790", x"f78d", x"f78a", x"f787", x"f784", x"f781", x"f77d", x"f77a", 
    x"f777", x"f774", x"f771", x"f76e", x"f76b", x"f767", x"f764", x"f761", 
    x"f75e", x"f75b", x"f758", x"f755", x"f752", x"f74e", x"f74b", x"f748", 
    x"f745", x"f742", x"f73f", x"f73c", x"f738", x"f735", x"f732", x"f72f", 
    x"f72c", x"f729", x"f726", x"f723", x"f71f", x"f71c", x"f719", x"f716", 
    x"f713", x"f710", x"f70d", x"f709", x"f706", x"f703", x"f700", x"f6fd", 
    x"f6fa", x"f6f7", x"f6f4", x"f6f0", x"f6ed", x"f6ea", x"f6e7", x"f6e4", 
    x"f6e1", x"f6de", x"f6da", x"f6d7", x"f6d4", x"f6d1", x"f6ce", x"f6cb", 
    x"f6c8", x"f6c5", x"f6c1", x"f6be", x"f6bb", x"f6b8", x"f6b5", x"f6b2", 
    x"f6af", x"f6ab", x"f6a8", x"f6a5", x"f6a2", x"f69f", x"f69c", x"f699", 
    x"f696", x"f692", x"f68f", x"f68c", x"f689", x"f686", x"f683", x"f680", 
    x"f67c", x"f679", x"f676", x"f673", x"f670", x"f66d", x"f66a", x"f667", 
    x"f663", x"f660", x"f65d", x"f65a", x"f657", x"f654", x"f651", x"f64d", 
    x"f64a", x"f647", x"f644", x"f641", x"f63e", x"f63b", x"f638", x"f634", 
    x"f631", x"f62e", x"f62b", x"f628", x"f625", x"f622", x"f61e", x"f61b", 
    x"f618", x"f615", x"f612", x"f60f", x"f60c", x"f609", x"f605", x"f602", 
    x"f5ff", x"f5fc", x"f5f9", x"f5f6", x"f5f3", x"f5ef", x"f5ec", x"f5e9", 
    x"f5e6", x"f5e3", x"f5e0", x"f5dd", x"f5da", x"f5d6", x"f5d3", x"f5d0", 
    x"f5cd", x"f5ca", x"f5c7", x"f5c4", x"f5c1", x"f5bd", x"f5ba", x"f5b7", 
    x"f5b4", x"f5b1", x"f5ae", x"f5ab", x"f5a7", x"f5a4", x"f5a1", x"f59e", 
    x"f59b", x"f598", x"f595", x"f592", x"f58e", x"f58b", x"f588", x"f585", 
    x"f582", x"f57f", x"f57c", x"f579", x"f575", x"f572", x"f56f", x"f56c", 
    x"f569", x"f566", x"f563", x"f55f", x"f55c", x"f559", x"f556", x"f553", 
    x"f550", x"f54d", x"f54a", x"f546", x"f543", x"f540", x"f53d", x"f53a", 
    x"f537", x"f534", x"f531", x"f52d", x"f52a", x"f527", x"f524", x"f521", 
    x"f51e", x"f51b", x"f517", x"f514", x"f511", x"f50e", x"f50b", x"f508", 
    x"f505", x"f502", x"f4fe", x"f4fb", x"f4f8", x"f4f5", x"f4f2", x"f4ef", 
    x"f4ec", x"f4e9", x"f4e5", x"f4e2", x"f4df", x"f4dc", x"f4d9", x"f4d6", 
    x"f4d3", x"f4cf", x"f4cc", x"f4c9", x"f4c6", x"f4c3", x"f4c0", x"f4bd", 
    x"f4ba", x"f4b6", x"f4b3", x"f4b0", x"f4ad", x"f4aa", x"f4a7", x"f4a4", 
    x"f4a1", x"f49d", x"f49a", x"f497", x"f494", x"f491", x"f48e", x"f48b", 
    x"f488", x"f484", x"f481", x"f47e", x"f47b", x"f478", x"f475", x"f472", 
    x"f46e", x"f46b", x"f468", x"f465", x"f462", x"f45f", x"f45c", x"f459", 
    x"f455", x"f452", x"f44f", x"f44c", x"f449", x"f446", x"f443", x"f440", 
    x"f43c", x"f439", x"f436", x"f433", x"f430", x"f42d", x"f42a", x"f427", 
    x"f423", x"f420", x"f41d", x"f41a", x"f417", x"f414", x"f411", x"f40d", 
    x"f40a", x"f407", x"f404", x"f401", x"f3fe", x"f3fb", x"f3f8", x"f3f4", 
    x"f3f1", x"f3ee", x"f3eb", x"f3e8", x"f3e5", x"f3e2", x"f3df", x"f3db", 
    x"f3d8", x"f3d5", x"f3d2", x"f3cf", x"f3cc", x"f3c9", x"f3c6", x"f3c2", 
    x"f3bf", x"f3bc", x"f3b9", x"f3b6", x"f3b3", x"f3b0", x"f3ad", x"f3a9", 
    x"f3a6", x"f3a3", x"f3a0", x"f39d", x"f39a", x"f397", x"f394", x"f390", 
    x"f38d", x"f38a", x"f387", x"f384", x"f381", x"f37e", x"f37b", x"f377", 
    x"f374", x"f371", x"f36e", x"f36b", x"f368", x"f365", x"f362", x"f35e", 
    x"f35b", x"f358", x"f355", x"f352", x"f34f", x"f34c", x"f349", x"f345", 
    x"f342", x"f33f", x"f33c", x"f339", x"f336", x"f333", x"f32f", x"f32c", 
    x"f329", x"f326", x"f323", x"f320", x"f31d", x"f31a", x"f316", x"f313", 
    x"f310", x"f30d", x"f30a", x"f307", x"f304", x"f301", x"f2fd", x"f2fa", 
    x"f2f7", x"f2f4", x"f2f1", x"f2ee", x"f2eb", x"f2e8", x"f2e4", x"f2e1", 
    x"f2de", x"f2db", x"f2d8", x"f2d5", x"f2d2", x"f2cf", x"f2cb", x"f2c8", 
    x"f2c5", x"f2c2", x"f2bf", x"f2bc", x"f2b9", x"f2b6", x"f2b2", x"f2af", 
    x"f2ac", x"f2a9", x"f2a6", x"f2a3", x"f2a0", x"f29d", x"f29a", x"f296", 
    x"f293", x"f290", x"f28d", x"f28a", x"f287", x"f284", x"f281", x"f27d", 
    x"f27a", x"f277", x"f274", x"f271", x"f26e", x"f26b", x"f268", x"f264", 
    x"f261", x"f25e", x"f25b", x"f258", x"f255", x"f252", x"f24f", x"f24b", 
    x"f248", x"f245", x"f242", x"f23f", x"f23c", x"f239", x"f236", x"f232", 
    x"f22f", x"f22c", x"f229", x"f226", x"f223", x"f220", x"f21d", x"f219", 
    x"f216", x"f213", x"f210", x"f20d", x"f20a", x"f207", x"f204", x"f200", 
    x"f1fd", x"f1fa", x"f1f7", x"f1f4", x"f1f1", x"f1ee", x"f1eb", x"f1e7", 
    x"f1e4", x"f1e1", x"f1de", x"f1db", x"f1d8", x"f1d5", x"f1d2", x"f1ce", 
    x"f1cb", x"f1c8", x"f1c5", x"f1c2", x"f1bf", x"f1bc", x"f1b9", x"f1b6", 
    x"f1b2", x"f1af", x"f1ac", x"f1a9", x"f1a6", x"f1a3", x"f1a0", x"f19d", 
    x"f199", x"f196", x"f193", x"f190", x"f18d", x"f18a", x"f187", x"f184", 
    x"f180", x"f17d", x"f17a", x"f177", x"f174", x"f171", x"f16e", x"f16b", 
    x"f167", x"f164", x"f161", x"f15e", x"f15b", x"f158", x"f155", x"f152", 
    x"f14f", x"f14b", x"f148", x"f145", x"f142", x"f13f", x"f13c", x"f139", 
    x"f136", x"f132", x"f12f", x"f12c", x"f129", x"f126", x"f123", x"f120", 
    x"f11d", x"f119", x"f116", x"f113", x"f110", x"f10d", x"f10a", x"f107", 
    x"f104", x"f101", x"f0fd", x"f0fa", x"f0f7", x"f0f4", x"f0f1", x"f0ee", 
    x"f0eb", x"f0e8", x"f0e4", x"f0e1", x"f0de", x"f0db", x"f0d8", x"f0d5", 
    x"f0d2", x"f0cf", x"f0cb", x"f0c8", x"f0c5", x"f0c2", x"f0bf", x"f0bc", 
    x"f0b9", x"f0b6", x"f0b3", x"f0af", x"f0ac", x"f0a9", x"f0a6", x"f0a3", 
    x"f0a0", x"f09d", x"f09a", x"f096", x"f093", x"f090", x"f08d", x"f08a", 
    x"f087", x"f084", x"f081", x"f07e", x"f07a", x"f077", x"f074", x"f071", 
    x"f06e", x"f06b", x"f068", x"f065", x"f061", x"f05e", x"f05b", x"f058", 
    x"f055", x"f052", x"f04f", x"f04c", x"f048", x"f045", x"f042", x"f03f", 
    x"f03c", x"f039", x"f036", x"f033", x"f030", x"f02c", x"f029", x"f026", 
    x"f023", x"f020", x"f01d", x"f01a", x"f017", x"f014", x"f010", x"f00d", 
    x"f00a", x"f007", x"f004", x"f001", x"effe", x"effb", x"eff7", x"eff4", 
    x"eff1", x"efee", x"efeb", x"efe8", x"efe5", x"efe2", x"efdf", x"efdb", 
    x"efd8", x"efd5", x"efd2", x"efcf", x"efcc", x"efc9", x"efc6", x"efc2", 
    x"efbf", x"efbc", x"efb9", x"efb6", x"efb3", x"efb0", x"efad", x"efaa", 
    x"efa6", x"efa3", x"efa0", x"ef9d", x"ef9a", x"ef97", x"ef94", x"ef91", 
    x"ef8e", x"ef8a", x"ef87", x"ef84", x"ef81", x"ef7e", x"ef7b", x"ef78", 
    x"ef75", x"ef71", x"ef6e", x"ef6b", x"ef68", x"ef65", x"ef62", x"ef5f", 
    x"ef5c", x"ef59", x"ef55", x"ef52", x"ef4f", x"ef4c", x"ef49", x"ef46", 
    x"ef43", x"ef40", x"ef3d", x"ef39", x"ef36", x"ef33", x"ef30", x"ef2d", 
    x"ef2a", x"ef27", x"ef24", x"ef20", x"ef1d", x"ef1a", x"ef17", x"ef14", 
    x"ef11", x"ef0e", x"ef0b", x"ef08", x"ef04", x"ef01", x"eefe", x"eefb", 
    x"eef8", x"eef5", x"eef2", x"eeef", x"eeec", x"eee8", x"eee5", x"eee2", 
    x"eedf", x"eedc", x"eed9", x"eed6", x"eed3", x"eed0", x"eecc", x"eec9", 
    x"eec6", x"eec3", x"eec0", x"eebd", x"eeba", x"eeb7", x"eeb4", x"eeb0", 
    x"eead", x"eeaa", x"eea7", x"eea4", x"eea1", x"ee9e", x"ee9b", x"ee98", 
    x"ee94", x"ee91", x"ee8e", x"ee8b", x"ee88", x"ee85", x"ee82", x"ee7f", 
    x"ee7b", x"ee78", x"ee75", x"ee72", x"ee6f", x"ee6c", x"ee69", x"ee66", 
    x"ee63", x"ee5f", x"ee5c", x"ee59", x"ee56", x"ee53", x"ee50", x"ee4d", 
    x"ee4a", x"ee47", x"ee43", x"ee40", x"ee3d", x"ee3a", x"ee37", x"ee34", 
    x"ee31", x"ee2e", x"ee2b", x"ee27", x"ee24", x"ee21", x"ee1e", x"ee1b", 
    x"ee18", x"ee15", x"ee12", x"ee0f", x"ee0b", x"ee08", x"ee05", x"ee02", 
    x"edff", x"edfc", x"edf9", x"edf6", x"edf3", x"edf0", x"edec", x"ede9", 
    x"ede6", x"ede3", x"ede0", x"eddd", x"edda", x"edd7", x"edd4", x"edd0", 
    x"edcd", x"edca", x"edc7", x"edc4", x"edc1", x"edbe", x"edbb", x"edb8", 
    x"edb4", x"edb1", x"edae", x"edab", x"eda8", x"eda5", x"eda2", x"ed9f", 
    x"ed9c", x"ed98", x"ed95", x"ed92", x"ed8f", x"ed8c", x"ed89", x"ed86", 
    x"ed83", x"ed80", x"ed7c", x"ed79", x"ed76", x"ed73", x"ed70", x"ed6d", 
    x"ed6a", x"ed67", x"ed64", x"ed60", x"ed5d", x"ed5a", x"ed57", x"ed54", 
    x"ed51", x"ed4e", x"ed4b", x"ed48", x"ed45", x"ed41", x"ed3e", x"ed3b", 
    x"ed38", x"ed35", x"ed32", x"ed2f", x"ed2c", x"ed29", x"ed25", x"ed22", 
    x"ed1f", x"ed1c", x"ed19", x"ed16", x"ed13", x"ed10", x"ed0d", x"ed09", 
    x"ed06", x"ed03", x"ed00", x"ecfd", x"ecfa", x"ecf7", x"ecf4", x"ecf1", 
    x"ecee", x"ecea", x"ece7", x"ece4", x"ece1", x"ecde", x"ecdb", x"ecd8", 
    x"ecd5", x"ecd2", x"ecce", x"eccb", x"ecc8", x"ecc5", x"ecc2", x"ecbf", 
    x"ecbc", x"ecb9", x"ecb6", x"ecb3", x"ecaf", x"ecac", x"eca9", x"eca6", 
    x"eca3", x"eca0", x"ec9d", x"ec9a", x"ec97", x"ec93", x"ec90", x"ec8d", 
    x"ec8a", x"ec87", x"ec84", x"ec81", x"ec7e", x"ec7b", x"ec78", x"ec74", 
    x"ec71", x"ec6e", x"ec6b", x"ec68", x"ec65", x"ec62", x"ec5f", x"ec5c", 
    x"ec58", x"ec55", x"ec52", x"ec4f", x"ec4c", x"ec49", x"ec46", x"ec43", 
    x"ec40", x"ec3d", x"ec39", x"ec36", x"ec33", x"ec30", x"ec2d", x"ec2a", 
    x"ec27", x"ec24", x"ec21", x"ec1d", x"ec1a", x"ec17", x"ec14", x"ec11", 
    x"ec0e", x"ec0b", x"ec08", x"ec05", x"ec02", x"ebfe", x"ebfb", x"ebf8", 
    x"ebf5", x"ebf2", x"ebef", x"ebec", x"ebe9", x"ebe6", x"ebe3", x"ebdf", 
    x"ebdc", x"ebd9", x"ebd6", x"ebd3", x"ebd0", x"ebcd", x"ebca", x"ebc7", 
    x"ebc4", x"ebc0", x"ebbd", x"ebba", x"ebb7", x"ebb4", x"ebb1", x"ebae", 
    x"ebab", x"eba8", x"eba4", x"eba1", x"eb9e", x"eb9b", x"eb98", x"eb95", 
    x"eb92", x"eb8f", x"eb8c", x"eb89", x"eb85", x"eb82", x"eb7f", x"eb7c", 
    x"eb79", x"eb76", x"eb73", x"eb70", x"eb6d", x"eb6a", x"eb66", x"eb63", 
    x"eb60", x"eb5d", x"eb5a", x"eb57", x"eb54", x"eb51", x"eb4e", x"eb4b", 
    x"eb47", x"eb44", x"eb41", x"eb3e", x"eb3b", x"eb38", x"eb35", x"eb32", 
    x"eb2f", x"eb2c", x"eb28", x"eb25", x"eb22", x"eb1f", x"eb1c", x"eb19", 
    x"eb16", x"eb13", x"eb10", x"eb0d", x"eb09", x"eb06", x"eb03", x"eb00", 
    x"eafd", x"eafa", x"eaf7", x"eaf4", x"eaf1", x"eaee", x"eaea", x"eae7", 
    x"eae4", x"eae1", x"eade", x"eadb", x"ead8", x"ead5", x"ead2", x"eacf", 
    x"eacc", x"eac8", x"eac5", x"eac2", x"eabf", x"eabc", x"eab9", x"eab6", 
    x"eab3", x"eab0", x"eaad", x"eaa9", x"eaa6", x"eaa3", x"eaa0", x"ea9d", 
    x"ea9a", x"ea97", x"ea94", x"ea91", x"ea8e", x"ea8a", x"ea87", x"ea84", 
    x"ea81", x"ea7e", x"ea7b", x"ea78", x"ea75", x"ea72", x"ea6f", x"ea6b", 
    x"ea68", x"ea65", x"ea62", x"ea5f", x"ea5c", x"ea59", x"ea56", x"ea53", 
    x"ea50", x"ea4d", x"ea49", x"ea46", x"ea43", x"ea40", x"ea3d", x"ea3a", 
    x"ea37", x"ea34", x"ea31", x"ea2e", x"ea2a", x"ea27", x"ea24", x"ea21", 
    x"ea1e", x"ea1b", x"ea18", x"ea15", x"ea12", x"ea0f", x"ea0c", x"ea08", 
    x"ea05", x"ea02", x"e9ff", x"e9fc", x"e9f9", x"e9f6", x"e9f3", x"e9f0", 
    x"e9ed", x"e9e9", x"e9e6", x"e9e3", x"e9e0", x"e9dd", x"e9da", x"e9d7", 
    x"e9d4", x"e9d1", x"e9ce", x"e9cb", x"e9c7", x"e9c4", x"e9c1", x"e9be", 
    x"e9bb", x"e9b8", x"e9b5", x"e9b2", x"e9af", x"e9ac", x"e9a9", x"e9a5", 
    x"e9a2", x"e99f", x"e99c", x"e999", x"e996", x"e993", x"e990", x"e98d", 
    x"e98a", x"e986", x"e983", x"e980", x"e97d", x"e97a", x"e977", x"e974", 
    x"e971", x"e96e", x"e96b", x"e968", x"e964", x"e961", x"e95e", x"e95b", 
    x"e958", x"e955", x"e952", x"e94f", x"e94c", x"e949", x"e946", x"e942", 
    x"e93f", x"e93c", x"e939", x"e936", x"e933", x"e930", x"e92d", x"e92a", 
    x"e927", x"e924", x"e920", x"e91d", x"e91a", x"e917", x"e914", x"e911", 
    x"e90e", x"e90b", x"e908", x"e905", x"e902", x"e8fe", x"e8fb", x"e8f8", 
    x"e8f5", x"e8f2", x"e8ef", x"e8ec", x"e8e9", x"e8e6", x"e8e3", x"e8e0", 
    x"e8dc", x"e8d9", x"e8d6", x"e8d3", x"e8d0", x"e8cd", x"e8ca", x"e8c7", 
    x"e8c4", x"e8c1", x"e8be", x"e8ba", x"e8b7", x"e8b4", x"e8b1", x"e8ae", 
    x"e8ab", x"e8a8", x"e8a5", x"e8a2", x"e89f", x"e89c", x"e899", x"e895", 
    x"e892", x"e88f", x"e88c", x"e889", x"e886", x"e883", x"e880", x"e87d", 
    x"e87a", x"e877", x"e873", x"e870", x"e86d", x"e86a", x"e867", x"e864", 
    x"e861", x"e85e", x"e85b", x"e858", x"e855", x"e851", x"e84e", x"e84b", 
    x"e848", x"e845", x"e842", x"e83f", x"e83c", x"e839", x"e836", x"e833", 
    x"e830", x"e82c", x"e829", x"e826", x"e823", x"e820", x"e81d", x"e81a", 
    x"e817", x"e814", x"e811", x"e80e", x"e80a", x"e807", x"e804", x"e801", 
    x"e7fe", x"e7fb", x"e7f8", x"e7f5", x"e7f2", x"e7ef", x"e7ec", x"e7e9", 
    x"e7e5", x"e7e2", x"e7df", x"e7dc", x"e7d9", x"e7d6", x"e7d3", x"e7d0", 
    x"e7cd", x"e7ca", x"e7c7", x"e7c4", x"e7c0", x"e7bd", x"e7ba", x"e7b7", 
    x"e7b4", x"e7b1", x"e7ae", x"e7ab", x"e7a8", x"e7a5", x"e7a2", x"e79f", 
    x"e79b", x"e798", x"e795", x"e792", x"e78f", x"e78c", x"e789", x"e786", 
    x"e783", x"e780", x"e77d", x"e77a", x"e776", x"e773", x"e770", x"e76d", 
    x"e76a", x"e767", x"e764", x"e761", x"e75e", x"e75b", x"e758", x"e755", 
    x"e751", x"e74e", x"e74b", x"e748", x"e745", x"e742", x"e73f", x"e73c", 
    x"e739", x"e736", x"e733", x"e730", x"e72c", x"e729", x"e726", x"e723", 
    x"e720", x"e71d", x"e71a", x"e717", x"e714", x"e711", x"e70e", x"e70b", 
    x"e707", x"e704", x"e701", x"e6fe", x"e6fb", x"e6f8", x"e6f5", x"e6f2", 
    x"e6ef", x"e6ec", x"e6e9", x"e6e6", x"e6e3", x"e6df", x"e6dc", x"e6d9", 
    x"e6d6", x"e6d3", x"e6d0", x"e6cd", x"e6ca", x"e6c7", x"e6c4", x"e6c1", 
    x"e6be", x"e6ba", x"e6b7", x"e6b4", x"e6b1", x"e6ae", x"e6ab", x"e6a8", 
    x"e6a5", x"e6a2", x"e69f", x"e69c", x"e699", x"e696", x"e692", x"e68f", 
    x"e68c", x"e689", x"e686", x"e683", x"e680", x"e67d", x"e67a", x"e677", 
    x"e674", x"e671", x"e66d", x"e66a", x"e667", x"e664", x"e661", x"e65e", 
    x"e65b", x"e658", x"e655", x"e652", x"e64f", x"e64c", x"e649", x"e645", 
    x"e642", x"e63f", x"e63c", x"e639", x"e636", x"e633", x"e630", x"e62d", 
    x"e62a", x"e627", x"e624", x"e621", x"e61d", x"e61a", x"e617", x"e614", 
    x"e611", x"e60e", x"e60b", x"e608", x"e605", x"e602", x"e5ff", x"e5fc", 
    x"e5f9", x"e5f5", x"e5f2", x"e5ef", x"e5ec", x"e5e9", x"e5e6", x"e5e3", 
    x"e5e0", x"e5dd", x"e5da", x"e5d7", x"e5d4", x"e5d1", x"e5ce", x"e5ca", 
    x"e5c7", x"e5c4", x"e5c1", x"e5be", x"e5bb", x"e5b8", x"e5b5", x"e5b2", 
    x"e5af", x"e5ac", x"e5a9", x"e5a6", x"e5a2", x"e59f", x"e59c", x"e599", 
    x"e596", x"e593", x"e590", x"e58d", x"e58a", x"e587", x"e584", x"e581", 
    x"e57e", x"e57b", x"e577", x"e574", x"e571", x"e56e", x"e56b", x"e568", 
    x"e565", x"e562", x"e55f", x"e55c", x"e559", x"e556", x"e553", x"e54f", 
    x"e54c", x"e549", x"e546", x"e543", x"e540", x"e53d", x"e53a", x"e537", 
    x"e534", x"e531", x"e52e", x"e52b", x"e528", x"e524", x"e521", x"e51e", 
    x"e51b", x"e518", x"e515", x"e512", x"e50f", x"e50c", x"e509", x"e506", 
    x"e503", x"e500", x"e4fd", x"e4f9", x"e4f6", x"e4f3", x"e4f0", x"e4ed", 
    x"e4ea", x"e4e7", x"e4e4", x"e4e1", x"e4de", x"e4db", x"e4d8", x"e4d5", 
    x"e4d2", x"e4cf", x"e4cb", x"e4c8", x"e4c5", x"e4c2", x"e4bf", x"e4bc", 
    x"e4b9", x"e4b6", x"e4b3", x"e4b0", x"e4ad", x"e4aa", x"e4a7", x"e4a4", 
    x"e4a0", x"e49d", x"e49a", x"e497", x"e494", x"e491", x"e48e", x"e48b", 
    x"e488", x"e485", x"e482", x"e47f", x"e47c", x"e479", x"e476", x"e472", 
    x"e46f", x"e46c", x"e469", x"e466", x"e463", x"e460", x"e45d", x"e45a", 
    x"e457", x"e454", x"e451", x"e44e", x"e44b", x"e447", x"e444", x"e441", 
    x"e43e", x"e43b", x"e438", x"e435", x"e432", x"e42f", x"e42c", x"e429", 
    x"e426", x"e423", x"e420", x"e41d", x"e419", x"e416", x"e413", x"e410", 
    x"e40d", x"e40a", x"e407", x"e404", x"e401", x"e3fe", x"e3fb", x"e3f8", 
    x"e3f5", x"e3f2", x"e3ef", x"e3ec", x"e3e8", x"e3e5", x"e3e2", x"e3df", 
    x"e3dc", x"e3d9", x"e3d6", x"e3d3", x"e3d0", x"e3cd", x"e3ca", x"e3c7", 
    x"e3c4", x"e3c1", x"e3be", x"e3ba", x"e3b7", x"e3b4", x"e3b1", x"e3ae", 
    x"e3ab", x"e3a8", x"e3a5", x"e3a2", x"e39f", x"e39c", x"e399", x"e396", 
    x"e393", x"e390", x"e38d", x"e389", x"e386", x"e383", x"e380", x"e37d", 
    x"e37a", x"e377", x"e374", x"e371", x"e36e", x"e36b", x"e368", x"e365", 
    x"e362", x"e35f", x"e35c", x"e358", x"e355", x"e352", x"e34f", x"e34c", 
    x"e349", x"e346", x"e343", x"e340", x"e33d", x"e33a", x"e337", x"e334", 
    x"e331", x"e32e", x"e32b", x"e327", x"e324", x"e321", x"e31e", x"e31b", 
    x"e318", x"e315", x"e312", x"e30f", x"e30c", x"e309", x"e306", x"e303", 
    x"e300", x"e2fd", x"e2fa", x"e2f7", x"e2f3", x"e2f0", x"e2ed", x"e2ea", 
    x"e2e7", x"e2e4", x"e2e1", x"e2de", x"e2db", x"e2d8", x"e2d5", x"e2d2", 
    x"e2cf", x"e2cc", x"e2c9", x"e2c6", x"e2c3", x"e2bf", x"e2bc", x"e2b9", 
    x"e2b6", x"e2b3", x"e2b0", x"e2ad", x"e2aa", x"e2a7", x"e2a4", x"e2a1", 
    x"e29e", x"e29b", x"e298", x"e295", x"e292", x"e28f", x"e28b", x"e288", 
    x"e285", x"e282", x"e27f", x"e27c", x"e279", x"e276", x"e273", x"e270", 
    x"e26d", x"e26a", x"e267", x"e264", x"e261", x"e25e", x"e25b", x"e258", 
    x"e254", x"e251", x"e24e", x"e24b", x"e248", x"e245", x"e242", x"e23f", 
    x"e23c", x"e239", x"e236", x"e233", x"e230", x"e22d", x"e22a", x"e227", 
    x"e224", x"e221", x"e21d", x"e21a", x"e217", x"e214", x"e211", x"e20e", 
    x"e20b", x"e208", x"e205", x"e202", x"e1ff", x"e1fc", x"e1f9", x"e1f6", 
    x"e1f3", x"e1f0", x"e1ed", x"e1ea", x"e1e7", x"e1e3", x"e1e0", x"e1dd", 
    x"e1da", x"e1d7", x"e1d4", x"e1d1", x"e1ce", x"e1cb", x"e1c8", x"e1c5", 
    x"e1c2", x"e1bf", x"e1bc", x"e1b9", x"e1b6", x"e1b3", x"e1b0", x"e1ac", 
    x"e1a9", x"e1a6", x"e1a3", x"e1a0", x"e19d", x"e19a", x"e197", x"e194", 
    x"e191", x"e18e", x"e18b", x"e188", x"e185", x"e182", x"e17f", x"e17c", 
    x"e179", x"e176", x"e173", x"e16f", x"e16c", x"e169", x"e166", x"e163", 
    x"e160", x"e15d", x"e15a", x"e157", x"e154", x"e151", x"e14e", x"e14b", 
    x"e148", x"e145", x"e142", x"e13f", x"e13c", x"e139", x"e136", x"e132", 
    x"e12f", x"e12c", x"e129", x"e126", x"e123", x"e120", x"e11d", x"e11a", 
    x"e117", x"e114", x"e111", x"e10e", x"e10b", x"e108", x"e105", x"e102", 
    x"e0ff", x"e0fc", x"e0f9", x"e0f6", x"e0f2", x"e0ef", x"e0ec", x"e0e9", 
    x"e0e6", x"e0e3", x"e0e0", x"e0dd", x"e0da", x"e0d7", x"e0d4", x"e0d1", 
    x"e0ce", x"e0cb", x"e0c8", x"e0c5", x"e0c2", x"e0bf", x"e0bc", x"e0b9", 
    x"e0b6", x"e0b2", x"e0af", x"e0ac", x"e0a9", x"e0a6", x"e0a3", x"e0a0", 
    x"e09d", x"e09a", x"e097", x"e094", x"e091", x"e08e", x"e08b", x"e088", 
    x"e085", x"e082", x"e07f", x"e07c", x"e079", x"e076", x"e073", x"e06f", 
    x"e06c", x"e069", x"e066", x"e063", x"e060", x"e05d", x"e05a", x"e057", 
    x"e054", x"e051", x"e04e", x"e04b", x"e048", x"e045", x"e042", x"e03f", 
    x"e03c", x"e039", x"e036", x"e033", x"e030", x"e02d", x"e029", x"e026", 
    x"e023", x"e020", x"e01d", x"e01a", x"e017", x"e014", x"e011", x"e00e", 
    x"e00b", x"e008", x"e005", x"e002", x"dfff", x"dffc", x"dff9", x"dff6", 
    x"dff3", x"dff0", x"dfed", x"dfea", x"dfe7", x"dfe4", x"dfe0", x"dfdd", 
    x"dfda", x"dfd7", x"dfd4", x"dfd1", x"dfce", x"dfcb", x"dfc8", x"dfc5", 
    x"dfc2", x"dfbf", x"dfbc", x"dfb9", x"dfb6", x"dfb3", x"dfb0", x"dfad", 
    x"dfaa", x"dfa7", x"dfa4", x"dfa1", x"df9e", x"df9b", x"df98", x"df94", 
    x"df91", x"df8e", x"df8b", x"df88", x"df85", x"df82", x"df7f", x"df7c", 
    x"df79", x"df76", x"df73", x"df70", x"df6d", x"df6a", x"df67", x"df64", 
    x"df61", x"df5e", x"df5b", x"df58", x"df55", x"df52", x"df4f", x"df4c", 
    x"df49", x"df45", x"df42", x"df3f", x"df3c", x"df39", x"df36", x"df33", 
    x"df30", x"df2d", x"df2a", x"df27", x"df24", x"df21", x"df1e", x"df1b", 
    x"df18", x"df15", x"df12", x"df0f", x"df0c", x"df09", x"df06", x"df03", 
    x"df00", x"defd", x"defa", x"def7", x"def4", x"def0", x"deed", x"deea", 
    x"dee7", x"dee4", x"dee1", x"dede", x"dedb", x"ded8", x"ded5", x"ded2", 
    x"decf", x"decc", x"dec9", x"dec6", x"dec3", x"dec0", x"debd", x"deba", 
    x"deb7", x"deb4", x"deb1", x"deae", x"deab", x"dea8", x"dea5", x"dea2", 
    x"de9f", x"de9c", x"de98", x"de95", x"de92", x"de8f", x"de8c", x"de89", 
    x"de86", x"de83", x"de80", x"de7d", x"de7a", x"de77", x"de74", x"de71", 
    x"de6e", x"de6b", x"de68", x"de65", x"de62", x"de5f", x"de5c", x"de59", 
    x"de56", x"de53", x"de50", x"de4d", x"de4a", x"de47", x"de44", x"de41", 
    x"de3e", x"de3b", x"de37", x"de34", x"de31", x"de2e", x"de2b", x"de28", 
    x"de25", x"de22", x"de1f", x"de1c", x"de19", x"de16", x"de13", x"de10", 
    x"de0d", x"de0a", x"de07", x"de04", x"de01", x"ddfe", x"ddfb", x"ddf8", 
    x"ddf5", x"ddf2", x"ddef", x"ddec", x"dde9", x"dde6", x"dde3", x"dde0", 
    x"dddd", x"ddda", x"ddd7", x"ddd4", x"ddd1", x"ddcd", x"ddca", x"ddc7", 
    x"ddc4", x"ddc1", x"ddbe", x"ddbb", x"ddb8", x"ddb5", x"ddb2", x"ddaf", 
    x"ddac", x"dda9", x"dda6", x"dda3", x"dda0", x"dd9d", x"dd9a", x"dd97", 
    x"dd94", x"dd91", x"dd8e", x"dd8b", x"dd88", x"dd85", x"dd82", x"dd7f", 
    x"dd7c", x"dd79", x"dd76", x"dd73", x"dd70", x"dd6d", x"dd6a", x"dd67", 
    x"dd64", x"dd61", x"dd5e", x"dd5b", x"dd57", x"dd54", x"dd51", x"dd4e", 
    x"dd4b", x"dd48", x"dd45", x"dd42", x"dd3f", x"dd3c", x"dd39", x"dd36", 
    x"dd33", x"dd30", x"dd2d", x"dd2a", x"dd27", x"dd24", x"dd21", x"dd1e", 
    x"dd1b", x"dd18", x"dd15", x"dd12", x"dd0f", x"dd0c", x"dd09", x"dd06", 
    x"dd03", x"dd00", x"dcfd", x"dcfa", x"dcf7", x"dcf4", x"dcf1", x"dcee", 
    x"dceb", x"dce8", x"dce5", x"dce2", x"dcdf", x"dcdc", x"dcd9", x"dcd6", 
    x"dcd2", x"dccf", x"dccc", x"dcc9", x"dcc6", x"dcc3", x"dcc0", x"dcbd", 
    x"dcba", x"dcb7", x"dcb4", x"dcb1", x"dcae", x"dcab", x"dca8", x"dca5", 
    x"dca2", x"dc9f", x"dc9c", x"dc99", x"dc96", x"dc93", x"dc90", x"dc8d", 
    x"dc8a", x"dc87", x"dc84", x"dc81", x"dc7e", x"dc7b", x"dc78", x"dc75", 
    x"dc72", x"dc6f", x"dc6c", x"dc69", x"dc66", x"dc63", x"dc60", x"dc5d", 
    x"dc5a", x"dc57", x"dc54", x"dc51", x"dc4e", x"dc4b", x"dc48", x"dc45", 
    x"dc42", x"dc3f", x"dc3c", x"dc39", x"dc36", x"dc33", x"dc30", x"dc2c", 
    x"dc29", x"dc26", x"dc23", x"dc20", x"dc1d", x"dc1a", x"dc17", x"dc14", 
    x"dc11", x"dc0e", x"dc0b", x"dc08", x"dc05", x"dc02", x"dbff", x"dbfc", 
    x"dbf9", x"dbf6", x"dbf3", x"dbf0", x"dbed", x"dbea", x"dbe7", x"dbe4", 
    x"dbe1", x"dbde", x"dbdb", x"dbd8", x"dbd5", x"dbd2", x"dbcf", x"dbcc", 
    x"dbc9", x"dbc6", x"dbc3", x"dbc0", x"dbbd", x"dbba", x"dbb7", x"dbb4", 
    x"dbb1", x"dbae", x"dbab", x"dba8", x"dba5", x"dba2", x"db9f", x"db9c", 
    x"db99", x"db96", x"db93", x"db90", x"db8d", x"db8a", x"db87", x"db84", 
    x"db81", x"db7e", x"db7b", x"db78", x"db75", x"db72", x"db6f", x"db6c", 
    x"db69", x"db66", x"db63", x"db60", x"db5d", x"db5a", x"db57", x"db54", 
    x"db51", x"db4e", x"db4b", x"db48", x"db45", x"db42", x"db3f", x"db3b", 
    x"db38", x"db35", x"db32", x"db2f", x"db2c", x"db29", x"db26", x"db23", 
    x"db20", x"db1d", x"db1a", x"db17", x"db14", x"db11", x"db0e", x"db0b", 
    x"db08", x"db05", x"db02", x"daff", x"dafc", x"daf9", x"daf6", x"daf3", 
    x"daf0", x"daed", x"daea", x"dae7", x"dae4", x"dae1", x"dade", x"dadb", 
    x"dad8", x"dad5", x"dad2", x"dacf", x"dacc", x"dac9", x"dac6", x"dac3", 
    x"dac0", x"dabd", x"daba", x"dab7", x"dab4", x"dab1", x"daae", x"daab", 
    x"daa8", x"daa5", x"daa2", x"da9f", x"da9c", x"da99", x"da96", x"da93", 
    x"da90", x"da8d", x"da8a", x"da87", x"da84", x"da81", x"da7e", x"da7b", 
    x"da78", x"da75", x"da72", x"da6f", x"da6c", x"da69", x"da66", x"da63", 
    x"da60", x"da5d", x"da5a", x"da57", x"da54", x"da51", x"da4e", x"da4b", 
    x"da48", x"da45", x"da42", x"da3f", x"da3c", x"da39", x"da36", x"da33", 
    x"da30", x"da2d", x"da2a", x"da27", x"da24", x"da21", x"da1e", x"da1b", 
    x"da18", x"da15", x"da12", x"da0f", x"da0c", x"da09", x"da06", x"da03", 
    x"da00", x"d9fd", x"d9fa", x"d9f7", x"d9f4", x"d9f1", x"d9ee", x"d9eb", 
    x"d9e8", x"d9e5", x"d9e2", x"d9df", x"d9dc", x"d9d9", x"d9d6", x"d9d3", 
    x"d9d0", x"d9cd", x"d9ca", x"d9c7", x"d9c4", x"d9c1", x"d9be", x"d9bb", 
    x"d9b8", x"d9b5", x"d9b2", x"d9af", x"d9ac", x"d9a9", x"d9a6", x"d9a3", 
    x"d9a0", x"d99d", x"d99a", x"d997", x"d994", x"d991", x"d98e", x"d98b", 
    x"d988", x"d985", x"d982", x"d97f", x"d97c", x"d979", x"d976", x"d973", 
    x"d970", x"d96d", x"d96a", x"d967", x"d964", x"d961", x"d95e", x"d95b", 
    x"d958", x"d955", x"d952", x"d94f", x"d94c", x"d949", x"d946", x"d943", 
    x"d940", x"d93d", x"d93a", x"d937", x"d934", x"d931", x"d92e", x"d92b", 
    x"d928", x"d925", x"d922", x"d91f", x"d91c", x"d919", x"d916", x"d913", 
    x"d910", x"d90d", x"d90a", x"d907", x"d904", x"d901", x"d8fe", x"d8fb", 
    x"d8f8", x"d8f5", x"d8f2", x"d8ef", x"d8ec", x"d8e9", x"d8e6", x"d8e3", 
    x"d8e0", x"d8dd", x"d8da", x"d8d7", x"d8d4", x"d8d1", x"d8cf", x"d8cc", 
    x"d8c9", x"d8c6", x"d8c3", x"d8c0", x"d8bd", x"d8ba", x"d8b7", x"d8b4", 
    x"d8b1", x"d8ae", x"d8ab", x"d8a8", x"d8a5", x"d8a2", x"d89f", x"d89c", 
    x"d899", x"d896", x"d893", x"d890", x"d88d", x"d88a", x"d887", x"d884", 
    x"d881", x"d87e", x"d87b", x"d878", x"d875", x"d872", x"d86f", x"d86c", 
    x"d869", x"d866", x"d863", x"d860", x"d85d", x"d85a", x"d857", x"d854", 
    x"d851", x"d84e", x"d84b", x"d848", x"d845", x"d842", x"d83f", x"d83c", 
    x"d839", x"d836", x"d833", x"d830", x"d82d", x"d82a", x"d827", x"d824", 
    x"d821", x"d81e", x"d81b", x"d818", x"d815", x"d812", x"d80f", x"d80c", 
    x"d809", x"d806", x"d803", x"d800", x"d7fd", x"d7fa", x"d7f7", x"d7f4", 
    x"d7f1", x"d7ee", x"d7eb", x"d7e9", x"d7e6", x"d7e3", x"d7e0", x"d7dd", 
    x"d7da", x"d7d7", x"d7d4", x"d7d1", x"d7ce", x"d7cb", x"d7c8", x"d7c5", 
    x"d7c2", x"d7bf", x"d7bc", x"d7b9", x"d7b6", x"d7b3", x"d7b0", x"d7ad", 
    x"d7aa", x"d7a7", x"d7a4", x"d7a1", x"d79e", x"d79b", x"d798", x"d795", 
    x"d792", x"d78f", x"d78c", x"d789", x"d786", x"d783", x"d780", x"d77d", 
    x"d77a", x"d777", x"d774", x"d771", x"d76e", x"d76b", x"d768", x"d765", 
    x"d762", x"d75f", x"d75c", x"d759", x"d756", x"d753", x"d750", x"d74d", 
    x"d74b", x"d748", x"d745", x"d742", x"d73f", x"d73c", x"d739", x"d736", 
    x"d733", x"d730", x"d72d", x"d72a", x"d727", x"d724", x"d721", x"d71e", 
    x"d71b", x"d718", x"d715", x"d712", x"d70f", x"d70c", x"d709", x"d706", 
    x"d703", x"d700", x"d6fd", x"d6fa", x"d6f7", x"d6f4", x"d6f1", x"d6ee", 
    x"d6eb", x"d6e8", x"d6e5", x"d6e2", x"d6df", x"d6dc", x"d6d9", x"d6d6", 
    x"d6d3", x"d6d0", x"d6ce", x"d6cb", x"d6c8", x"d6c5", x"d6c2", x"d6bf", 
    x"d6bc", x"d6b9", x"d6b6", x"d6b3", x"d6b0", x"d6ad", x"d6aa", x"d6a7", 
    x"d6a4", x"d6a1", x"d69e", x"d69b", x"d698", x"d695", x"d692", x"d68f", 
    x"d68c", x"d689", x"d686", x"d683", x"d680", x"d67d", x"d67a", x"d677", 
    x"d674", x"d671", x"d66e", x"d66b", x"d668", x"d665", x"d662", x"d660", 
    x"d65d", x"d65a", x"d657", x"d654", x"d651", x"d64e", x"d64b", x"d648", 
    x"d645", x"d642", x"d63f", x"d63c", x"d639", x"d636", x"d633", x"d630", 
    x"d62d", x"d62a", x"d627", x"d624", x"d621", x"d61e", x"d61b", x"d618", 
    x"d615", x"d612", x"d60f", x"d60c", x"d609", x"d606", x"d603", x"d601", 
    x"d5fe", x"d5fb", x"d5f8", x"d5f5", x"d5f2", x"d5ef", x"d5ec", x"d5e9", 
    x"d5e6", x"d5e3", x"d5e0", x"d5dd", x"d5da", x"d5d7", x"d5d4", x"d5d1", 
    x"d5ce", x"d5cb", x"d5c8", x"d5c5", x"d5c2", x"d5bf", x"d5bc", x"d5b9", 
    x"d5b6", x"d5b3", x"d5b0", x"d5ad", x"d5aa", x"d5a8", x"d5a5", x"d5a2", 
    x"d59f", x"d59c", x"d599", x"d596", x"d593", x"d590", x"d58d", x"d58a", 
    x"d587", x"d584", x"d581", x"d57e", x"d57b", x"d578", x"d575", x"d572", 
    x"d56f", x"d56c", x"d569", x"d566", x"d563", x"d560", x"d55d", x"d55a", 
    x"d558", x"d555", x"d552", x"d54f", x"d54c", x"d549", x"d546", x"d543", 
    x"d540", x"d53d", x"d53a", x"d537", x"d534", x"d531", x"d52e", x"d52b", 
    x"d528", x"d525", x"d522", x"d51f", x"d51c", x"d519", x"d516", x"d513", 
    x"d510", x"d50e", x"d50b", x"d508", x"d505", x"d502", x"d4ff", x"d4fc", 
    x"d4f9", x"d4f6", x"d4f3", x"d4f0", x"d4ed", x"d4ea", x"d4e7", x"d4e4", 
    x"d4e1", x"d4de", x"d4db", x"d4d8", x"d4d5", x"d4d2", x"d4cf", x"d4cc", 
    x"d4c9", x"d4c7", x"d4c4", x"d4c1", x"d4be", x"d4bb", x"d4b8", x"d4b5", 
    x"d4b2", x"d4af", x"d4ac", x"d4a9", x"d4a6", x"d4a3", x"d4a0", x"d49d", 
    x"d49a", x"d497", x"d494", x"d491", x"d48e", x"d48b", x"d488", x"d485", 
    x"d483", x"d480", x"d47d", x"d47a", x"d477", x"d474", x"d471", x"d46e", 
    x"d46b", x"d468", x"d465", x"d462", x"d45f", x"d45c", x"d459", x"d456", 
    x"d453", x"d450", x"d44d", x"d44a", x"d447", x"d445", x"d442", x"d43f", 
    x"d43c", x"d439", x"d436", x"d433", x"d430", x"d42d", x"d42a", x"d427", 
    x"d424", x"d421", x"d41e", x"d41b", x"d418", x"d415", x"d412", x"d40f", 
    x"d40c", x"d409", x"d407", x"d404", x"d401", x"d3fe", x"d3fb", x"d3f8", 
    x"d3f5", x"d3f2", x"d3ef", x"d3ec", x"d3e9", x"d3e6", x"d3e3", x"d3e0", 
    x"d3dd", x"d3da", x"d3d7", x"d3d4", x"d3d1", x"d3ce", x"d3cc", x"d3c9", 
    x"d3c6", x"d3c3", x"d3c0", x"d3bd", x"d3ba", x"d3b7", x"d3b4", x"d3b1", 
    x"d3ae", x"d3ab", x"d3a8", x"d3a5", x"d3a2", x"d39f", x"d39c", x"d399", 
    x"d396", x"d394", x"d391", x"d38e", x"d38b", x"d388", x"d385", x"d382", 
    x"d37f", x"d37c", x"d379", x"d376", x"d373", x"d370", x"d36d", x"d36a", 
    x"d367", x"d364", x"d361", x"d35f", x"d35c", x"d359", x"d356", x"d353", 
    x"d350", x"d34d", x"d34a", x"d347", x"d344", x"d341", x"d33e", x"d33b", 
    x"d338", x"d335", x"d332", x"d32f", x"d32c", x"d32a", x"d327", x"d324", 
    x"d321", x"d31e", x"d31b", x"d318", x"d315", x"d312", x"d30f", x"d30c", 
    x"d309", x"d306", x"d303", x"d300", x"d2fd", x"d2fa", x"d2f8", x"d2f5", 
    x"d2f2", x"d2ef", x"d2ec", x"d2e9", x"d2e6", x"d2e3", x"d2e0", x"d2dd", 
    x"d2da", x"d2d7", x"d2d4", x"d2d1", x"d2ce", x"d2cb", x"d2c9", x"d2c6", 
    x"d2c3", x"d2c0", x"d2bd", x"d2ba", x"d2b7", x"d2b4", x"d2b1", x"d2ae", 
    x"d2ab", x"d2a8", x"d2a5", x"d2a2", x"d29f", x"d29c", x"d299", x"d297", 
    x"d294", x"d291", x"d28e", x"d28b", x"d288", x"d285", x"d282", x"d27f", 
    x"d27c", x"d279", x"d276", x"d273", x"d270", x"d26d", x"d26b", x"d268", 
    x"d265", x"d262", x"d25f", x"d25c", x"d259", x"d256", x"d253", x"d250", 
    x"d24d", x"d24a", x"d247", x"d244", x"d241", x"d23e", x"d23c", x"d239", 
    x"d236", x"d233", x"d230", x"d22d", x"d22a", x"d227", x"d224", x"d221", 
    x"d21e", x"d21b", x"d218", x"d215", x"d212", x"d210", x"d20d", x"d20a", 
    x"d207", x"d204", x"d201", x"d1fe", x"d1fb", x"d1f8", x"d1f5", x"d1f2", 
    x"d1ef", x"d1ec", x"d1e9", x"d1e7", x"d1e4", x"d1e1", x"d1de", x"d1db", 
    x"d1d8", x"d1d5", x"d1d2", x"d1cf", x"d1cc", x"d1c9", x"d1c6", x"d1c3", 
    x"d1c0", x"d1be", x"d1bb", x"d1b8", x"d1b5", x"d1b2", x"d1af", x"d1ac", 
    x"d1a9", x"d1a6", x"d1a3", x"d1a0", x"d19d", x"d19a", x"d197", x"d195", 
    x"d192", x"d18f", x"d18c", x"d189", x"d186", x"d183", x"d180", x"d17d", 
    x"d17a", x"d177", x"d174", x"d171", x"d16e", x"d16c", x"d169", x"d166", 
    x"d163", x"d160", x"d15d", x"d15a", x"d157", x"d154", x"d151", x"d14e", 
    x"d14b", x"d148", x"d146", x"d143", x"d140", x"d13d", x"d13a", x"d137", 
    x"d134", x"d131", x"d12e", x"d12b", x"d128", x"d125", x"d122", x"d11f", 
    x"d11d", x"d11a", x"d117", x"d114", x"d111", x"d10e", x"d10b", x"d108", 
    x"d105", x"d102", x"d0ff", x"d0fc", x"d0fa", x"d0f7", x"d0f4", x"d0f1", 
    x"d0ee", x"d0eb", x"d0e8", x"d0e5", x"d0e2", x"d0df", x"d0dc", x"d0d9", 
    x"d0d6", x"d0d4", x"d0d1", x"d0ce", x"d0cb", x"d0c8", x"d0c5", x"d0c2", 
    x"d0bf", x"d0bc", x"d0b9", x"d0b6", x"d0b3", x"d0b0", x"d0ae", x"d0ab", 
    x"d0a8", x"d0a5", x"d0a2", x"d09f", x"d09c", x"d099", x"d096", x"d093", 
    x"d090", x"d08d", x"d08b", x"d088", x"d085", x"d082", x"d07f", x"d07c", 
    x"d079", x"d076", x"d073", x"d070", x"d06d", x"d06a", x"d068", x"d065", 
    x"d062", x"d05f", x"d05c", x"d059", x"d056", x"d053", x"d050", x"d04d", 
    x"d04a", x"d047", x"d045", x"d042", x"d03f", x"d03c", x"d039", x"d036", 
    x"d033", x"d030", x"d02d", x"d02a", x"d027", x"d025", x"d022", x"d01f", 
    x"d01c", x"d019", x"d016", x"d013", x"d010", x"d00d", x"d00a", x"d007", 
    x"d004", x"d002", x"cfff", x"cffc", x"cff9", x"cff6", x"cff3", x"cff0", 
    x"cfed", x"cfea", x"cfe7", x"cfe4", x"cfe2", x"cfdf", x"cfdc", x"cfd9", 
    x"cfd6", x"cfd3", x"cfd0", x"cfcd", x"cfca", x"cfc7", x"cfc4", x"cfc2", 
    x"cfbf", x"cfbc", x"cfb9", x"cfb6", x"cfb3", x"cfb0", x"cfad", x"cfaa", 
    x"cfa7", x"cfa4", x"cfa2", x"cf9f", x"cf9c", x"cf99", x"cf96", x"cf93", 
    x"cf90", x"cf8d", x"cf8a", x"cf87", x"cf84", x"cf82", x"cf7f", x"cf7c", 
    x"cf79", x"cf76", x"cf73", x"cf70", x"cf6d", x"cf6a", x"cf67", x"cf64", 
    x"cf62", x"cf5f", x"cf5c", x"cf59", x"cf56", x"cf53", x"cf50", x"cf4d", 
    x"cf4a", x"cf47", x"cf44", x"cf42", x"cf3f", x"cf3c", x"cf39", x"cf36", 
    x"cf33", x"cf30", x"cf2d", x"cf2a", x"cf27", x"cf25", x"cf22", x"cf1f", 
    x"cf1c", x"cf19", x"cf16", x"cf13", x"cf10", x"cf0d", x"cf0a", x"cf08", 
    x"cf05", x"cf02", x"ceff", x"cefc", x"cef9", x"cef6", x"cef3", x"cef0", 
    x"ceed", x"ceea", x"cee8", x"cee5", x"cee2", x"cedf", x"cedc", x"ced9", 
    x"ced6", x"ced3", x"ced0", x"cecd", x"cecb", x"cec8", x"cec5", x"cec2", 
    x"cebf", x"cebc", x"ceb9", x"ceb6", x"ceb3", x"ceb0", x"ceae", x"ceab", 
    x"cea8", x"cea5", x"cea2", x"ce9f", x"ce9c", x"ce99", x"ce96", x"ce94", 
    x"ce91", x"ce8e", x"ce8b", x"ce88", x"ce85", x"ce82", x"ce7f", x"ce7c", 
    x"ce79", x"ce77", x"ce74", x"ce71", x"ce6e", x"ce6b", x"ce68", x"ce65", 
    x"ce62", x"ce5f", x"ce5c", x"ce5a", x"ce57", x"ce54", x"ce51", x"ce4e", 
    x"ce4b", x"ce48", x"ce45", x"ce42", x"ce40", x"ce3d", x"ce3a", x"ce37", 
    x"ce34", x"ce31", x"ce2e", x"ce2b", x"ce28", x"ce25", x"ce23", x"ce20", 
    x"ce1d", x"ce1a", x"ce17", x"ce14", x"ce11", x"ce0e", x"ce0b", x"ce09", 
    x"ce06", x"ce03", x"ce00", x"cdfd", x"cdfa", x"cdf7", x"cdf4", x"cdf1", 
    x"cdef", x"cdec", x"cde9", x"cde6", x"cde3", x"cde0", x"cddd", x"cdda", 
    x"cdd7", x"cdd5", x"cdd2", x"cdcf", x"cdcc", x"cdc9", x"cdc6", x"cdc3", 
    x"cdc0", x"cdbd", x"cdba", x"cdb8", x"cdb5", x"cdb2", x"cdaf", x"cdac", 
    x"cda9", x"cda6", x"cda3", x"cda1", x"cd9e", x"cd9b", x"cd98", x"cd95", 
    x"cd92", x"cd8f", x"cd8c", x"cd89", x"cd87", x"cd84", x"cd81", x"cd7e", 
    x"cd7b", x"cd78", x"cd75", x"cd72", x"cd6f", x"cd6d", x"cd6a", x"cd67", 
    x"cd64", x"cd61", x"cd5e", x"cd5b", x"cd58", x"cd55", x"cd53", x"cd50", 
    x"cd4d", x"cd4a", x"cd47", x"cd44", x"cd41", x"cd3e", x"cd3b", x"cd39", 
    x"cd36", x"cd33", x"cd30", x"cd2d", x"cd2a", x"cd27", x"cd24", x"cd22", 
    x"cd1f", x"cd1c", x"cd19", x"cd16", x"cd13", x"cd10", x"cd0d", x"cd0a", 
    x"cd08", x"cd05", x"cd02", x"ccff", x"ccfc", x"ccf9", x"ccf6", x"ccf3", 
    x"ccf1", x"ccee", x"cceb", x"cce8", x"cce5", x"cce2", x"ccdf", x"ccdc", 
    x"ccda", x"ccd7", x"ccd4", x"ccd1", x"ccce", x"cccb", x"ccc8", x"ccc5", 
    x"ccc2", x"ccc0", x"ccbd", x"ccba", x"ccb7", x"ccb4", x"ccb1", x"ccae", 
    x"ccab", x"cca9", x"cca6", x"cca3", x"cca0", x"cc9d", x"cc9a", x"cc97", 
    x"cc94", x"cc92", x"cc8f", x"cc8c", x"cc89", x"cc86", x"cc83", x"cc80", 
    x"cc7d", x"cc7b", x"cc78", x"cc75", x"cc72", x"cc6f", x"cc6c", x"cc69", 
    x"cc66", x"cc64", x"cc61", x"cc5e", x"cc5b", x"cc58", x"cc55", x"cc52", 
    x"cc4f", x"cc4d", x"cc4a", x"cc47", x"cc44", x"cc41", x"cc3e", x"cc3b", 
    x"cc38", x"cc36", x"cc33", x"cc30", x"cc2d", x"cc2a", x"cc27", x"cc24", 
    x"cc21", x"cc1f", x"cc1c", x"cc19", x"cc16", x"cc13", x"cc10", x"cc0d", 
    x"cc0a", x"cc08", x"cc05", x"cc02", x"cbff", x"cbfc", x"cbf9", x"cbf6", 
    x"cbf4", x"cbf1", x"cbee", x"cbeb", x"cbe8", x"cbe5", x"cbe2", x"cbdf", 
    x"cbdd", x"cbda", x"cbd7", x"cbd4", x"cbd1", x"cbce", x"cbcb", x"cbc8", 
    x"cbc6", x"cbc3", x"cbc0", x"cbbd", x"cbba", x"cbb7", x"cbb4", x"cbb2", 
    x"cbaf", x"cbac", x"cba9", x"cba6", x"cba3", x"cba0", x"cb9d", x"cb9b", 
    x"cb98", x"cb95", x"cb92", x"cb8f", x"cb8c", x"cb89", x"cb87", x"cb84", 
    x"cb81", x"cb7e", x"cb7b", x"cb78", x"cb75", x"cb72", x"cb70", x"cb6d", 
    x"cb6a", x"cb67", x"cb64", x"cb61", x"cb5e", x"cb5c", x"cb59", x"cb56", 
    x"cb53", x"cb50", x"cb4d", x"cb4a", x"cb48", x"cb45", x"cb42", x"cb3f", 
    x"cb3c", x"cb39", x"cb36", x"cb34", x"cb31", x"cb2e", x"cb2b", x"cb28", 
    x"cb25", x"cb22", x"cb1f", x"cb1d", x"cb1a", x"cb17", x"cb14", x"cb11", 
    x"cb0e", x"cb0b", x"cb09", x"cb06", x"cb03", x"cb00", x"cafd", x"cafa", 
    x"caf7", x"caf5", x"caf2", x"caef", x"caec", x"cae9", x"cae6", x"cae3", 
    x"cae1", x"cade", x"cadb", x"cad8", x"cad5", x"cad2", x"cacf", x"cacd", 
    x"caca", x"cac7", x"cac4", x"cac1", x"cabe", x"cabb", x"cab9", x"cab6", 
    x"cab3", x"cab0", x"caad", x"caaa", x"caa7", x"caa5", x"caa2", x"ca9f", 
    x"ca9c", x"ca99", x"ca96", x"ca93", x"ca91", x"ca8e", x"ca8b", x"ca88", 
    x"ca85", x"ca82", x"ca7f", x"ca7d", x"ca7a", x"ca77", x"ca74", x"ca71", 
    x"ca6e", x"ca6b", x"ca69", x"ca66", x"ca63", x"ca60", x"ca5d", x"ca5a", 
    x"ca58", x"ca55", x"ca52", x"ca4f", x"ca4c", x"ca49", x"ca46", x"ca44", 
    x"ca41", x"ca3e", x"ca3b", x"ca38", x"ca35", x"ca32", x"ca30", x"ca2d", 
    x"ca2a", x"ca27", x"ca24", x"ca21", x"ca1f", x"ca1c", x"ca19", x"ca16", 
    x"ca13", x"ca10", x"ca0d", x"ca0b", x"ca08", x"ca05", x"ca02", x"c9ff", 
    x"c9fc", x"c9f9", x"c9f7", x"c9f4", x"c9f1", x"c9ee", x"c9eb", x"c9e8", 
    x"c9e6", x"c9e3", x"c9e0", x"c9dd", x"c9da", x"c9d7", x"c9d4", x"c9d2", 
    x"c9cf", x"c9cc", x"c9c9", x"c9c6", x"c9c3", x"c9c1", x"c9be", x"c9bb", 
    x"c9b8", x"c9b5", x"c9b2", x"c9af", x"c9ad", x"c9aa", x"c9a7", x"c9a4", 
    x"c9a1", x"c99e", x"c99c", x"c999", x"c996", x"c993", x"c990", x"c98d", 
    x"c98a", x"c988", x"c985", x"c982", x"c97f", x"c97c", x"c979", x"c977", 
    x"c974", x"c971", x"c96e", x"c96b", x"c968", x"c966", x"c963", x"c960", 
    x"c95d", x"c95a", x"c957", x"c955", x"c952", x"c94f", x"c94c", x"c949", 
    x"c946", x"c943", x"c941", x"c93e", x"c93b", x"c938", x"c935", x"c932", 
    x"c930", x"c92d", x"c92a", x"c927", x"c924", x"c921", x"c91f", x"c91c", 
    x"c919", x"c916", x"c913", x"c910", x"c90e", x"c90b", x"c908", x"c905", 
    x"c902", x"c8ff", x"c8fd", x"c8fa", x"c8f7", x"c8f4", x"c8f1", x"c8ee", 
    x"c8eb", x"c8e9", x"c8e6", x"c8e3", x"c8e0", x"c8dd", x"c8da", x"c8d8", 
    x"c8d5", x"c8d2", x"c8cf", x"c8cc", x"c8c9", x"c8c7", x"c8c4", x"c8c1", 
    x"c8be", x"c8bb", x"c8b8", x"c8b6", x"c8b3", x"c8b0", x"c8ad", x"c8aa", 
    x"c8a7", x"c8a5", x"c8a2", x"c89f", x"c89c", x"c899", x"c896", x"c894", 
    x"c891", x"c88e", x"c88b", x"c888", x"c885", x"c883", x"c880", x"c87d", 
    x"c87a", x"c877", x"c875", x"c872", x"c86f", x"c86c", x"c869", x"c866", 
    x"c864", x"c861", x"c85e", x"c85b", x"c858", x"c855", x"c853", x"c850", 
    x"c84d", x"c84a", x"c847", x"c844", x"c842", x"c83f", x"c83c", x"c839", 
    x"c836", x"c833", x"c831", x"c82e", x"c82b", x"c828", x"c825", x"c822", 
    x"c820", x"c81d", x"c81a", x"c817", x"c814", x"c812", x"c80f", x"c80c", 
    x"c809", x"c806", x"c803", x"c801", x"c7fe", x"c7fb", x"c7f8", x"c7f5", 
    x"c7f2", x"c7f0", x"c7ed", x"c7ea", x"c7e7", x"c7e4", x"c7e2", x"c7df", 
    x"c7dc", x"c7d9", x"c7d6", x"c7d3", x"c7d1", x"c7ce", x"c7cb", x"c7c8", 
    x"c7c5", x"c7c2", x"c7c0", x"c7bd", x"c7ba", x"c7b7", x"c7b4", x"c7b2", 
    x"c7af", x"c7ac", x"c7a9", x"c7a6", x"c7a3", x"c7a1", x"c79e", x"c79b", 
    x"c798", x"c795", x"c793", x"c790", x"c78d", x"c78a", x"c787", x"c784", 
    x"c782", x"c77f", x"c77c", x"c779", x"c776", x"c773", x"c771", x"c76e", 
    x"c76b", x"c768", x"c765", x"c763", x"c760", x"c75d", x"c75a", x"c757", 
    x"c755", x"c752", x"c74f", x"c74c", x"c749", x"c746", x"c744", x"c741", 
    x"c73e", x"c73b", x"c738", x"c736", x"c733", x"c730", x"c72d", x"c72a", 
    x"c727", x"c725", x"c722", x"c71f", x"c71c", x"c719", x"c717", x"c714", 
    x"c711", x"c70e", x"c70b", x"c708", x"c706", x"c703", x"c700", x"c6fd", 
    x"c6fa", x"c6f8", x"c6f5", x"c6f2", x"c6ef", x"c6ec", x"c6ea", x"c6e7", 
    x"c6e4", x"c6e1", x"c6de", x"c6dc", x"c6d9", x"c6d6", x"c6d3", x"c6d0", 
    x"c6cd", x"c6cb", x"c6c8", x"c6c5", x"c6c2", x"c6bf", x"c6bd", x"c6ba", 
    x"c6b7", x"c6b4", x"c6b1", x"c6af", x"c6ac", x"c6a9", x"c6a6", x"c6a3", 
    x"c6a0", x"c69e", x"c69b", x"c698", x"c695", x"c692", x"c690", x"c68d", 
    x"c68a", x"c687", x"c684", x"c682", x"c67f", x"c67c", x"c679", x"c676", 
    x"c674", x"c671", x"c66e", x"c66b", x"c668", x"c666", x"c663", x"c660", 
    x"c65d", x"c65a", x"c658", x"c655", x"c652", x"c64f", x"c64c", x"c64a", 
    x"c647", x"c644", x"c641", x"c63e", x"c63b", x"c639", x"c636", x"c633", 
    x"c630", x"c62d", x"c62b", x"c628", x"c625", x"c622", x"c61f", x"c61d", 
    x"c61a", x"c617", x"c614", x"c611", x"c60f", x"c60c", x"c609", x"c606", 
    x"c603", x"c601", x"c5fe", x"c5fb", x"c5f8", x"c5f5", x"c5f3", x"c5f0", 
    x"c5ed", x"c5ea", x"c5e7", x"c5e5", x"c5e2", x"c5df", x"c5dc", x"c5d9", 
    x"c5d7", x"c5d4", x"c5d1", x"c5ce", x"c5cb", x"c5c9", x"c5c6", x"c5c3", 
    x"c5c0", x"c5bd", x"c5bb", x"c5b8", x"c5b5", x"c5b2", x"c5af", x"c5ad", 
    x"c5aa", x"c5a7", x"c5a4", x"c5a2", x"c59f", x"c59c", x"c599", x"c596", 
    x"c594", x"c591", x"c58e", x"c58b", x"c588", x"c586", x"c583", x"c580", 
    x"c57d", x"c57a", x"c578", x"c575", x"c572", x"c56f", x"c56c", x"c56a", 
    x"c567", x"c564", x"c561", x"c55e", x"c55c", x"c559", x"c556", x"c553", 
    x"c550", x"c54e", x"c54b", x"c548", x"c545", x"c543", x"c540", x"c53d", 
    x"c53a", x"c537", x"c535", x"c532", x"c52f", x"c52c", x"c529", x"c527", 
    x"c524", x"c521", x"c51e", x"c51b", x"c519", x"c516", x"c513", x"c510", 
    x"c50e", x"c50b", x"c508", x"c505", x"c502", x"c500", x"c4fd", x"c4fa", 
    x"c4f7", x"c4f4", x"c4f2", x"c4ef", x"c4ec", x"c4e9", x"c4e7", x"c4e4", 
    x"c4e1", x"c4de", x"c4db", x"c4d9", x"c4d6", x"c4d3", x"c4d0", x"c4cd", 
    x"c4cb", x"c4c8", x"c4c5", x"c4c2", x"c4c0", x"c4bd", x"c4ba", x"c4b7", 
    x"c4b4", x"c4b2", x"c4af", x"c4ac", x"c4a9", x"c4a6", x"c4a4", x"c4a1", 
    x"c49e", x"c49b", x"c499", x"c496", x"c493", x"c490", x"c48d", x"c48b", 
    x"c488", x"c485", x"c482", x"c47f", x"c47d", x"c47a", x"c477", x"c474", 
    x"c472", x"c46f", x"c46c", x"c469", x"c466", x"c464", x"c461", x"c45e", 
    x"c45b", x"c459", x"c456", x"c453", x"c450", x"c44d", x"c44b", x"c448", 
    x"c445", x"c442", x"c440", x"c43d", x"c43a", x"c437", x"c434", x"c432", 
    x"c42f", x"c42c", x"c429", x"c427", x"c424", x"c421", x"c41e", x"c41b", 
    x"c419", x"c416", x"c413", x"c410", x"c40e", x"c40b", x"c408", x"c405", 
    x"c402", x"c400", x"c3fd", x"c3fa", x"c3f7", x"c3f5", x"c3f2", x"c3ef", 
    x"c3ec", x"c3ea", x"c3e7", x"c3e4", x"c3e1", x"c3de", x"c3dc", x"c3d9", 
    x"c3d6", x"c3d3", x"c3d1", x"c3ce", x"c3cb", x"c3c8", x"c3c5", x"c3c3", 
    x"c3c0", x"c3bd", x"c3ba", x"c3b8", x"c3b5", x"c3b2", x"c3af", x"c3ad", 
    x"c3aa", x"c3a7", x"c3a4", x"c3a1", x"c39f", x"c39c", x"c399", x"c396", 
    x"c394", x"c391", x"c38e", x"c38b", x"c389", x"c386", x"c383", x"c380", 
    x"c37d", x"c37b", x"c378", x"c375", x"c372", x"c370", x"c36d", x"c36a", 
    x"c367", x"c365", x"c362", x"c35f", x"c35c", x"c359", x"c357", x"c354", 
    x"c351", x"c34e", x"c34c", x"c349", x"c346", x"c343", x"c341", x"c33e", 
    x"c33b", x"c338", x"c336", x"c333", x"c330", x"c32d", x"c32a", x"c328", 
    x"c325", x"c322", x"c31f", x"c31d", x"c31a", x"c317", x"c314", x"c312", 
    x"c30f", x"c30c", x"c309", x"c307", x"c304", x"c301", x"c2fe", x"c2fb", 
    x"c2f9", x"c2f6", x"c2f3", x"c2f0", x"c2ee", x"c2eb", x"c2e8", x"c2e5", 
    x"c2e3", x"c2e0", x"c2dd", x"c2da", x"c2d8", x"c2d5", x"c2d2", x"c2cf", 
    x"c2cd", x"c2ca", x"c2c7", x"c2c4", x"c2c2", x"c2bf", x"c2bc", x"c2b9", 
    x"c2b6", x"c2b4", x"c2b1", x"c2ae", x"c2ab", x"c2a9", x"c2a6", x"c2a3", 
    x"c2a0", x"c29e", x"c29b", x"c298", x"c295", x"c293", x"c290", x"c28d", 
    x"c28a", x"c288", x"c285", x"c282", x"c27f", x"c27d", x"c27a", x"c277", 
    x"c274", x"c272", x"c26f", x"c26c", x"c269", x"c267", x"c264", x"c261", 
    x"c25e", x"c25c", x"c259", x"c256", x"c253", x"c251", x"c24e", x"c24b", 
    x"c248", x"c246", x"c243", x"c240", x"c23d", x"c23b", x"c238", x"c235", 
    x"c232", x"c230", x"c22d", x"c22a", x"c227", x"c225", x"c222", x"c21f", 
    x"c21c", x"c21a", x"c217", x"c214", x"c211", x"c20f", x"c20c", x"c209", 
    x"c206", x"c204", x"c201", x"c1fe", x"c1fb", x"c1f9", x"c1f6", x"c1f3", 
    x"c1f0", x"c1ee", x"c1eb", x"c1e8", x"c1e5", x"c1e3", x"c1e0", x"c1dd", 
    x"c1da", x"c1d8", x"c1d5", x"c1d2", x"c1cf", x"c1cd", x"c1ca", x"c1c7", 
    x"c1c4", x"c1c2", x"c1bf", x"c1bc", x"c1b9", x"c1b7", x"c1b4", x"c1b1", 
    x"c1ae", x"c1ac", x"c1a9", x"c1a6", x"c1a3", x"c1a1", x"c19e", x"c19b", 
    x"c198", x"c196", x"c193", x"c190", x"c18d", x"c18b", x"c188", x"c185", 
    x"c183", x"c180", x"c17d", x"c17a", x"c178", x"c175", x"c172", x"c16f", 
    x"c16d", x"c16a", x"c167", x"c164", x"c162", x"c15f", x"c15c", x"c159", 
    x"c157", x"c154", x"c151", x"c14e", x"c14c", x"c149", x"c146", x"c143", 
    x"c141", x"c13e", x"c13b", x"c139", x"c136", x"c133", x"c130", x"c12e", 
    x"c12b", x"c128", x"c125", x"c123", x"c120", x"c11d", x"c11a", x"c118", 
    x"c115", x"c112", x"c10f", x"c10d", x"c10a", x"c107", x"c105", x"c102", 
    x"c0ff", x"c0fc", x"c0fa", x"c0f7", x"c0f4", x"c0f1", x"c0ef", x"c0ec", 
    x"c0e9", x"c0e6", x"c0e4", x"c0e1", x"c0de", x"c0dc", x"c0d9", x"c0d6", 
    x"c0d3", x"c0d1", x"c0ce", x"c0cb", x"c0c8", x"c0c6", x"c0c3", x"c0c0", 
    x"c0bd", x"c0bb", x"c0b8", x"c0b5", x"c0b3", x"c0b0", x"c0ad", x"c0aa", 
    x"c0a8", x"c0a5", x"c0a2", x"c09f", x"c09d", x"c09a", x"c097", x"c095", 
    x"c092", x"c08f", x"c08c", x"c08a", x"c087", x"c084", x"c081", x"c07f", 
    x"c07c", x"c079", x"c077", x"c074", x"c071", x"c06e", x"c06c", x"c069", 
    x"c066", x"c063", x"c061", x"c05e", x"c05b", x"c059", x"c056", x"c053", 
    x"c050", x"c04e", x"c04b", x"c048", x"c045", x"c043", x"c040", x"c03d", 
    x"c03b", x"c038", x"c035", x"c032", x"c030", x"c02d", x"c02a", x"c028", 
    x"c025", x"c022", x"c01f", x"c01d", x"c01a", x"c017", x"c014", x"c012", 
    x"c00f", x"c00c", x"c00a", x"c007", x"c004", x"c001", x"bfff", x"bffc", 
    x"bff9", x"bff7", x"bff4", x"bff1", x"bfee", x"bfec", x"bfe9", x"bfe6", 
    x"bfe3", x"bfe1", x"bfde", x"bfdb", x"bfd9", x"bfd6", x"bfd3", x"bfd0", 
    x"bfce", x"bfcb", x"bfc8", x"bfc6", x"bfc3", x"bfc0", x"bfbd", x"bfbb", 
    x"bfb8", x"bfb5", x"bfb3", x"bfb0", x"bfad", x"bfaa", x"bfa8", x"bfa5", 
    x"bfa2", x"bfa0", x"bf9d", x"bf9a", x"bf97", x"bf95", x"bf92", x"bf8f", 
    x"bf8d", x"bf8a", x"bf87", x"bf84", x"bf82", x"bf7f", x"bf7c", x"bf7a", 
    x"bf77", x"bf74", x"bf71", x"bf6f", x"bf6c", x"bf69", x"bf67", x"bf64", 
    x"bf61", x"bf5e", x"bf5c", x"bf59", x"bf56", x"bf54", x"bf51", x"bf4e", 
    x"bf4b", x"bf49", x"bf46", x"bf43", x"bf41", x"bf3e", x"bf3b", x"bf38", 
    x"bf36", x"bf33", x"bf30", x"bf2e", x"bf2b", x"bf28", x"bf26", x"bf23", 
    x"bf20", x"bf1d", x"bf1b", x"bf18", x"bf15", x"bf13", x"bf10", x"bf0d", 
    x"bf0a", x"bf08", x"bf05", x"bf02", x"bf00", x"befd", x"befa", x"bef8", 
    x"bef5", x"bef2", x"beef", x"beed", x"beea", x"bee7", x"bee5", x"bee2", 
    x"bedf", x"bedc", x"beda", x"bed7", x"bed4", x"bed2", x"becf", x"becc", 
    x"beca", x"bec7", x"bec4", x"bec1", x"bebf", x"bebc", x"beb9", x"beb7", 
    x"beb4", x"beb1", x"beaf", x"beac", x"bea9", x"bea6", x"bea4", x"bea1", 
    x"be9e", x"be9c", x"be99", x"be96", x"be93", x"be91", x"be8e", x"be8b", 
    x"be89", x"be86", x"be83", x"be81", x"be7e", x"be7b", x"be79", x"be76", 
    x"be73", x"be70", x"be6e", x"be6b", x"be68", x"be66", x"be63", x"be60", 
    x"be5e", x"be5b", x"be58", x"be55", x"be53", x"be50", x"be4d", x"be4b", 
    x"be48", x"be45", x"be43", x"be40", x"be3d", x"be3a", x"be38", x"be35", 
    x"be32", x"be30", x"be2d", x"be2a", x"be28", x"be25", x"be22", x"be20", 
    x"be1d", x"be1a", x"be17", x"be15", x"be12", x"be0f", x"be0d", x"be0a", 
    x"be07", x"be05", x"be02", x"bdff", x"bdfd", x"bdfa", x"bdf7", x"bdf4", 
    x"bdf2", x"bdef", x"bdec", x"bdea", x"bde7", x"bde4", x"bde2", x"bddf", 
    x"bddc", x"bdda", x"bdd7", x"bdd4", x"bdd1", x"bdcf", x"bdcc", x"bdc9", 
    x"bdc7", x"bdc4", x"bdc1", x"bdbf", x"bdbc", x"bdb9", x"bdb7", x"bdb4", 
    x"bdb1", x"bdaf", x"bdac", x"bda9", x"bda6", x"bda4", x"bda1", x"bd9e", 
    x"bd9c", x"bd99", x"bd96", x"bd94", x"bd91", x"bd8e", x"bd8c", x"bd89", 
    x"bd86", x"bd84", x"bd81", x"bd7e", x"bd7c", x"bd79", x"bd76", x"bd73", 
    x"bd71", x"bd6e", x"bd6b", x"bd69", x"bd66", x"bd63", x"bd61", x"bd5e", 
    x"bd5b", x"bd59", x"bd56", x"bd53", x"bd51", x"bd4e", x"bd4b", x"bd49", 
    x"bd46", x"bd43", x"bd41", x"bd3e", x"bd3b", x"bd38", x"bd36", x"bd33", 
    x"bd30", x"bd2e", x"bd2b", x"bd28", x"bd26", x"bd23", x"bd20", x"bd1e", 
    x"bd1b", x"bd18", x"bd16", x"bd13", x"bd10", x"bd0e", x"bd0b", x"bd08", 
    x"bd06", x"bd03", x"bd00", x"bcfe", x"bcfb", x"bcf8", x"bcf6", x"bcf3", 
    x"bcf0", x"bced", x"bceb", x"bce8", x"bce5", x"bce3", x"bce0", x"bcdd", 
    x"bcdb", x"bcd8", x"bcd5", x"bcd3", x"bcd0", x"bccd", x"bccb", x"bcc8", 
    x"bcc5", x"bcc3", x"bcc0", x"bcbd", x"bcbb", x"bcb8", x"bcb5", x"bcb3", 
    x"bcb0", x"bcad", x"bcab", x"bca8", x"bca5", x"bca3", x"bca0", x"bc9d", 
    x"bc9b", x"bc98", x"bc95", x"bc93", x"bc90", x"bc8d", x"bc8b", x"bc88", 
    x"bc85", x"bc83", x"bc80", x"bc7d", x"bc7b", x"bc78", x"bc75", x"bc73", 
    x"bc70", x"bc6d", x"bc6b", x"bc68", x"bc65", x"bc63", x"bc60", x"bc5d", 
    x"bc5b", x"bc58", x"bc55", x"bc53", x"bc50", x"bc4d", x"bc4b", x"bc48", 
    x"bc45", x"bc43", x"bc40", x"bc3d", x"bc3b", x"bc38", x"bc35", x"bc33", 
    x"bc30", x"bc2d", x"bc2b", x"bc28", x"bc25", x"bc23", x"bc20", x"bc1d", 
    x"bc1b", x"bc18", x"bc15", x"bc13", x"bc10", x"bc0d", x"bc0b", x"bc08", 
    x"bc05", x"bc03", x"bc00", x"bbfd", x"bbfb", x"bbf8", x"bbf5", x"bbf3", 
    x"bbf0", x"bbed", x"bbeb", x"bbe8", x"bbe5", x"bbe3", x"bbe0", x"bbdd", 
    x"bbdb", x"bbd8", x"bbd5", x"bbd3", x"bbd0", x"bbcd", x"bbcb", x"bbc8", 
    x"bbc5", x"bbc3", x"bbc0", x"bbbe", x"bbbb", x"bbb8", x"bbb6", x"bbb3", 
    x"bbb0", x"bbae", x"bbab", x"bba8", x"bba6", x"bba3", x"bba0", x"bb9e", 
    x"bb9b", x"bb98", x"bb96", x"bb93", x"bb90", x"bb8e", x"bb8b", x"bb88", 
    x"bb86", x"bb83", x"bb80", x"bb7e", x"bb7b", x"bb78", x"bb76", x"bb73", 
    x"bb71", x"bb6e", x"bb6b", x"bb69", x"bb66", x"bb63", x"bb61", x"bb5e", 
    x"bb5b", x"bb59", x"bb56", x"bb53", x"bb51", x"bb4e", x"bb4b", x"bb49", 
    x"bb46", x"bb43", x"bb41", x"bb3e", x"bb3b", x"bb39", x"bb36", x"bb34", 
    x"bb31", x"bb2e", x"bb2c", x"bb29", x"bb26", x"bb24", x"bb21", x"bb1e", 
    x"bb1c", x"bb19", x"bb16", x"bb14", x"bb11", x"bb0e", x"bb0c", x"bb09", 
    x"bb07", x"bb04", x"bb01", x"baff", x"bafc", x"baf9", x"baf7", x"baf4", 
    x"baf1", x"baef", x"baec", x"bae9", x"bae7", x"bae4", x"bae1", x"badf", 
    x"badc", x"bada", x"bad7", x"bad4", x"bad2", x"bacf", x"bacc", x"baca", 
    x"bac7", x"bac4", x"bac2", x"babf", x"babc", x"baba", x"bab7", x"bab5", 
    x"bab2", x"baaf", x"baad", x"baaa", x"baa7", x"baa5", x"baa2", x"ba9f", 
    x"ba9d", x"ba9a", x"ba98", x"ba95", x"ba92", x"ba90", x"ba8d", x"ba8a", 
    x"ba88", x"ba85", x"ba82", x"ba80", x"ba7d", x"ba7a", x"ba78", x"ba75", 
    x"ba73", x"ba70", x"ba6d", x"ba6b", x"ba68", x"ba65", x"ba63", x"ba60", 
    x"ba5d", x"ba5b", x"ba58", x"ba56", x"ba53", x"ba50", x"ba4e", x"ba4b", 
    x"ba48", x"ba46", x"ba43", x"ba41", x"ba3e", x"ba3b", x"ba39", x"ba36", 
    x"ba33", x"ba31", x"ba2e", x"ba2b", x"ba29", x"ba26", x"ba24", x"ba21", 
    x"ba1e", x"ba1c", x"ba19", x"ba16", x"ba14", x"ba11", x"ba0e", x"ba0c", 
    x"ba09", x"ba07", x"ba04", x"ba01", x"b9ff", x"b9fc", x"b9f9", x"b9f7", 
    x"b9f4", x"b9f2", x"b9ef", x"b9ec", x"b9ea", x"b9e7", x"b9e4", x"b9e2", 
    x"b9df", x"b9dd", x"b9da", x"b9d7", x"b9d5", x"b9d2", x"b9cf", x"b9cd", 
    x"b9ca", x"b9c8", x"b9c5", x"b9c2", x"b9c0", x"b9bd", x"b9ba", x"b9b8", 
    x"b9b5", x"b9b3", x"b9b0", x"b9ad", x"b9ab", x"b9a8", x"b9a5", x"b9a3", 
    x"b9a0", x"b99e", x"b99b", x"b998", x"b996", x"b993", x"b990", x"b98e", 
    x"b98b", x"b989", x"b986", x"b983", x"b981", x"b97e", x"b97b", x"b979", 
    x"b976", x"b974", x"b971", x"b96e", x"b96c", x"b969", x"b966", x"b964", 
    x"b961", x"b95f", x"b95c", x"b959", x"b957", x"b954", x"b951", x"b94f", 
    x"b94c", x"b94a", x"b947", x"b944", x"b942", x"b93f", x"b93d", x"b93a", 
    x"b937", x"b935", x"b932", x"b92f", x"b92d", x"b92a", x"b928", x"b925", 
    x"b922", x"b920", x"b91d", x"b91b", x"b918", x"b915", x"b913", x"b910", 
    x"b90d", x"b90b", x"b908", x"b906", x"b903", x"b900", x"b8fe", x"b8fb", 
    x"b8f9", x"b8f6", x"b8f3", x"b8f1", x"b8ee", x"b8eb", x"b8e9", x"b8e6", 
    x"b8e4", x"b8e1", x"b8de", x"b8dc", x"b8d9", x"b8d7", x"b8d4", x"b8d1", 
    x"b8cf", x"b8cc", x"b8ca", x"b8c7", x"b8c4", x"b8c2", x"b8bf", x"b8bc", 
    x"b8ba", x"b8b7", x"b8b5", x"b8b2", x"b8af", x"b8ad", x"b8aa", x"b8a8", 
    x"b8a5", x"b8a2", x"b8a0", x"b89d", x"b89b", x"b898", x"b895", x"b893", 
    x"b890", x"b88e", x"b88b", x"b888", x"b886", x"b883", x"b880", x"b87e", 
    x"b87b", x"b879", x"b876", x"b873", x"b871", x"b86e", x"b86c", x"b869", 
    x"b866", x"b864", x"b861", x"b85f", x"b85c", x"b859", x"b857", x"b854", 
    x"b852", x"b84f", x"b84c", x"b84a", x"b847", x"b845", x"b842", x"b83f", 
    x"b83d", x"b83a", x"b838", x"b835", x"b832", x"b830", x"b82d", x"b82b", 
    x"b828", x"b825", x"b823", x"b820", x"b81e", x"b81b", x"b818", x"b816", 
    x"b813", x"b811", x"b80e", x"b80b", x"b809", x"b806", x"b804", x"b801", 
    x"b7fe", x"b7fc", x"b7f9", x"b7f7", x"b7f4", x"b7f1", x"b7ef", x"b7ec", 
    x"b7ea", x"b7e7", x"b7e4", x"b7e2", x"b7df", x"b7dd", x"b7da", x"b7d7", 
    x"b7d5", x"b7d2", x"b7d0", x"b7cd", x"b7cb", x"b7c8", x"b7c5", x"b7c3", 
    x"b7c0", x"b7be", x"b7bb", x"b7b8", x"b7b6", x"b7b3", x"b7b1", x"b7ae", 
    x"b7ab", x"b7a9", x"b7a6", x"b7a4", x"b7a1", x"b79e", x"b79c", x"b799", 
    x"b797", x"b794", x"b791", x"b78f", x"b78c", x"b78a", x"b787", x"b785", 
    x"b782", x"b77f", x"b77d", x"b77a", x"b778", x"b775", x"b772", x"b770", 
    x"b76d", x"b76b", x"b768", x"b765", x"b763", x"b760", x"b75e", x"b75b", 
    x"b759", x"b756", x"b753", x"b751", x"b74e", x"b74c", x"b749", x"b746", 
    x"b744", x"b741", x"b73f", x"b73c", x"b73a", x"b737", x"b734", x"b732", 
    x"b72f", x"b72d", x"b72a", x"b727", x"b725", x"b722", x"b720", x"b71d", 
    x"b71b", x"b718", x"b715", x"b713", x"b710", x"b70e", x"b70b", x"b708", 
    x"b706", x"b703", x"b701", x"b6fe", x"b6fc", x"b6f9", x"b6f6", x"b6f4", 
    x"b6f1", x"b6ef", x"b6ec", x"b6e9", x"b6e7", x"b6e4", x"b6e2", x"b6df", 
    x"b6dd", x"b6da", x"b6d7", x"b6d5", x"b6d2", x"b6d0", x"b6cd", x"b6cb", 
    x"b6c8", x"b6c5", x"b6c3", x"b6c0", x"b6be", x"b6bb", x"b6b9", x"b6b6", 
    x"b6b3", x"b6b1", x"b6ae", x"b6ac", x"b6a9", x"b6a6", x"b6a4", x"b6a1", 
    x"b69f", x"b69c", x"b69a", x"b697", x"b694", x"b692", x"b68f", x"b68d", 
    x"b68a", x"b688", x"b685", x"b682", x"b680", x"b67d", x"b67b", x"b678", 
    x"b676", x"b673", x"b670", x"b66e", x"b66b", x"b669", x"b666", x"b664", 
    x"b661", x"b65e", x"b65c", x"b659", x"b657", x"b654", x"b652", x"b64f", 
    x"b64c", x"b64a", x"b647", x"b645", x"b642", x"b640", x"b63d", x"b63b", 
    x"b638", x"b635", x"b633", x"b630", x"b62e", x"b62b", x"b629", x"b626", 
    x"b623", x"b621", x"b61e", x"b61c", x"b619", x"b617", x"b614", x"b611", 
    x"b60f", x"b60c", x"b60a", x"b607", x"b605", x"b602", x"b600", x"b5fd", 
    x"b5fa", x"b5f8", x"b5f5", x"b5f3", x"b5f0", x"b5ee", x"b5eb", x"b5e8", 
    x"b5e6", x"b5e3", x"b5e1", x"b5de", x"b5dc", x"b5d9", x"b5d7", x"b5d4", 
    x"b5d1", x"b5cf", x"b5cc", x"b5ca", x"b5c7", x"b5c5", x"b5c2", x"b5bf", 
    x"b5bd", x"b5ba", x"b5b8", x"b5b5", x"b5b3", x"b5b0", x"b5ae", x"b5ab", 
    x"b5a8", x"b5a6", x"b5a3", x"b5a1", x"b59e", x"b59c", x"b599", x"b597", 
    x"b594", x"b591", x"b58f", x"b58c", x"b58a", x"b587", x"b585", x"b582", 
    x"b580", x"b57d", x"b57a", x"b578", x"b575", x"b573", x"b570", x"b56e", 
    x"b56b", x"b569", x"b566", x"b563", x"b561", x"b55e", x"b55c", x"b559", 
    x"b557", x"b554", x"b552", x"b54f", x"b54d", x"b54a", x"b547", x"b545", 
    x"b542", x"b540", x"b53d", x"b53b", x"b538", x"b536", x"b533", x"b530", 
    x"b52e", x"b52b", x"b529", x"b526", x"b524", x"b521", x"b51f", x"b51c", 
    x"b51a", x"b517", x"b514", x"b512", x"b50f", x"b50d", x"b50a", x"b508", 
    x"b505", x"b503", x"b500", x"b4fe", x"b4fb", x"b4f8", x"b4f6", x"b4f3", 
    x"b4f1", x"b4ee", x"b4ec", x"b4e9", x"b4e7", x"b4e4", x"b4e2", x"b4df", 
    x"b4dc", x"b4da", x"b4d7", x"b4d5", x"b4d2", x"b4d0", x"b4cd", x"b4cb", 
    x"b4c8", x"b4c6", x"b4c3", x"b4c0", x"b4be", x"b4bb", x"b4b9", x"b4b6", 
    x"b4b4", x"b4b1", x"b4af", x"b4ac", x"b4aa", x"b4a7", x"b4a5", x"b4a2", 
    x"b49f", x"b49d", x"b49a", x"b498", x"b495", x"b493", x"b490", x"b48e", 
    x"b48b", x"b489", x"b486", x"b484", x"b481", x"b47e", x"b47c", x"b479", 
    x"b477", x"b474", x"b472", x"b46f", x"b46d", x"b46a", x"b468", x"b465", 
    x"b463", x"b460", x"b45e", x"b45b", x"b458", x"b456", x"b453", x"b451", 
    x"b44e", x"b44c", x"b449", x"b447", x"b444", x"b442", x"b43f", x"b43d", 
    x"b43a", x"b438", x"b435", x"b432", x"b430", x"b42d", x"b42b", x"b428", 
    x"b426", x"b423", x"b421", x"b41e", x"b41c", x"b419", x"b417", x"b414", 
    x"b412", x"b40f", x"b40c", x"b40a", x"b407", x"b405", x"b402", x"b400", 
    x"b3fd", x"b3fb", x"b3f8", x"b3f6", x"b3f3", x"b3f1", x"b3ee", x"b3ec", 
    x"b3e9", x"b3e7", x"b3e4", x"b3e2", x"b3df", x"b3dc", x"b3da", x"b3d7", 
    x"b3d5", x"b3d2", x"b3d0", x"b3cd", x"b3cb", x"b3c8", x"b3c6", x"b3c3", 
    x"b3c1", x"b3be", x"b3bc", x"b3b9", x"b3b7", x"b3b4", x"b3b2", x"b3af", 
    x"b3ad", x"b3aa", x"b3a7", x"b3a5", x"b3a2", x"b3a0", x"b39d", x"b39b", 
    x"b398", x"b396", x"b393", x"b391", x"b38e", x"b38c", x"b389", x"b387", 
    x"b384", x"b382", x"b37f", x"b37d", x"b37a", x"b378", x"b375", x"b373", 
    x"b370", x"b36e", x"b36b", x"b369", x"b366", x"b363", x"b361", x"b35e", 
    x"b35c", x"b359", x"b357", x"b354", x"b352", x"b34f", x"b34d", x"b34a", 
    x"b348", x"b345", x"b343", x"b340", x"b33e", x"b33b", x"b339", x"b336", 
    x"b334", x"b331", x"b32f", x"b32c", x"b32a", x"b327", x"b325", x"b322", 
    x"b320", x"b31d", x"b31b", x"b318", x"b316", x"b313", x"b311", x"b30e", 
    x"b30c", x"b309", x"b306", x"b304", x"b301", x"b2ff", x"b2fc", x"b2fa", 
    x"b2f7", x"b2f5", x"b2f2", x"b2f0", x"b2ed", x"b2eb", x"b2e8", x"b2e6", 
    x"b2e3", x"b2e1", x"b2de", x"b2dc", x"b2d9", x"b2d7", x"b2d4", x"b2d2", 
    x"b2cf", x"b2cd", x"b2ca", x"b2c8", x"b2c5", x"b2c3", x"b2c0", x"b2be", 
    x"b2bb", x"b2b9", x"b2b6", x"b2b4", x"b2b1", x"b2af", x"b2ac", x"b2aa", 
    x"b2a7", x"b2a5", x"b2a2", x"b2a0", x"b29d", x"b29b", x"b298", x"b296", 
    x"b293", x"b291", x"b28e", x"b28c", x"b289", x"b287", x"b284", x"b282", 
    x"b27f", x"b27d", x"b27a", x"b278", x"b275", x"b273", x"b270", x"b26e", 
    x"b26b", x"b269", x"b266", x"b264", x"b261", x"b25f", x"b25c", x"b25a", 
    x"b257", x"b255", x"b252", x"b250", x"b24d", x"b24b", x"b248", x"b246", 
    x"b243", x"b241", x"b23e", x"b23c", x"b239", x"b237", x"b234", x"b232", 
    x"b22f", x"b22d", x"b22a", x"b228", x"b225", x"b223", x"b220", x"b21e", 
    x"b21b", x"b219", x"b216", x"b214", x"b211", x"b20f", x"b20c", x"b20a", 
    x"b207", x"b205", x"b202", x"b200", x"b1fd", x"b1fb", x"b1f8", x"b1f6", 
    x"b1f3", x"b1f1", x"b1ef", x"b1ec", x"b1ea", x"b1e7", x"b1e5", x"b1e2", 
    x"b1e0", x"b1dd", x"b1db", x"b1d8", x"b1d6", x"b1d3", x"b1d1", x"b1ce", 
    x"b1cc", x"b1c9", x"b1c7", x"b1c4", x"b1c2", x"b1bf", x"b1bd", x"b1ba", 
    x"b1b8", x"b1b5", x"b1b3", x"b1b0", x"b1ae", x"b1ab", x"b1a9", x"b1a6", 
    x"b1a4", x"b1a1", x"b19f", x"b19c", x"b19a", x"b198", x"b195", x"b193", 
    x"b190", x"b18e", x"b18b", x"b189", x"b186", x"b184", x"b181", x"b17f", 
    x"b17c", x"b17a", x"b177", x"b175", x"b172", x"b170", x"b16d", x"b16b", 
    x"b168", x"b166", x"b163", x"b161", x"b15e", x"b15c", x"b159", x"b157", 
    x"b155", x"b152", x"b150", x"b14d", x"b14b", x"b148", x"b146", x"b143", 
    x"b141", x"b13e", x"b13c", x"b139", x"b137", x"b134", x"b132", x"b12f", 
    x"b12d", x"b12a", x"b128", x"b125", x"b123", x"b121", x"b11e", x"b11c", 
    x"b119", x"b117", x"b114", x"b112", x"b10f", x"b10d", x"b10a", x"b108", 
    x"b105", x"b103", x"b100", x"b0fe", x"b0fb", x"b0f9", x"b0f6", x"b0f4", 
    x"b0f2", x"b0ef", x"b0ed", x"b0ea", x"b0e8", x"b0e5", x"b0e3", x"b0e0", 
    x"b0de", x"b0db", x"b0d9", x"b0d6", x"b0d4", x"b0d1", x"b0cf", x"b0cd", 
    x"b0ca", x"b0c8", x"b0c5", x"b0c3", x"b0c0", x"b0be", x"b0bb", x"b0b9", 
    x"b0b6", x"b0b4", x"b0b1", x"b0af", x"b0ac", x"b0aa", x"b0a8", x"b0a5", 
    x"b0a3", x"b0a0", x"b09e", x"b09b", x"b099", x"b096", x"b094", x"b091", 
    x"b08f", x"b08c", x"b08a", x"b087", x"b085", x"b083", x"b080", x"b07e", 
    x"b07b", x"b079", x"b076", x"b074", x"b071", x"b06f", x"b06c", x"b06a", 
    x"b067", x"b065", x"b063", x"b060", x"b05e", x"b05b", x"b059", x"b056", 
    x"b054", x"b051", x"b04f", x"b04c", x"b04a", x"b048", x"b045", x"b043", 
    x"b040", x"b03e", x"b03b", x"b039", x"b036", x"b034", x"b031", x"b02f", 
    x"b02c", x"b02a", x"b028", x"b025", x"b023", x"b020", x"b01e", x"b01b", 
    x"b019", x"b016", x"b014", x"b011", x"b00f", x"b00d", x"b00a", x"b008", 
    x"b005", x"b003", x"b000", x"affe", x"affb", x"aff9", x"aff7", x"aff4", 
    x"aff2", x"afef", x"afed", x"afea", x"afe8", x"afe5", x"afe3", x"afe0", 
    x"afde", x"afdc", x"afd9", x"afd7", x"afd4", x"afd2", x"afcf", x"afcd", 
    x"afca", x"afc8", x"afc6", x"afc3", x"afc1", x"afbe", x"afbc", x"afb9", 
    x"afb7", x"afb4", x"afb2", x"afb0", x"afad", x"afab", x"afa8", x"afa6", 
    x"afa3", x"afa1", x"af9e", x"af9c", x"af99", x"af97", x"af95", x"af92", 
    x"af90", x"af8d", x"af8b", x"af88", x"af86", x"af84", x"af81", x"af7f", 
    x"af7c", x"af7a", x"af77", x"af75", x"af72", x"af70", x"af6e", x"af6b", 
    x"af69", x"af66", x"af64", x"af61", x"af5f", x"af5c", x"af5a", x"af58", 
    x"af55", x"af53", x"af50", x"af4e", x"af4b", x"af49", x"af46", x"af44", 
    x"af42", x"af3f", x"af3d", x"af3a", x"af38", x"af35", x"af33", x"af31", 
    x"af2e", x"af2c", x"af29", x"af27", x"af24", x"af22", x"af20", x"af1d", 
    x"af1b", x"af18", x"af16", x"af13", x"af11", x"af0e", x"af0c", x"af0a", 
    x"af07", x"af05", x"af02", x"af00", x"aefd", x"aefb", x"aef9", x"aef6", 
    x"aef4", x"aef1", x"aeef", x"aeec", x"aeea", x"aee8", x"aee5", x"aee3", 
    x"aee0", x"aede", x"aedb", x"aed9", x"aed7", x"aed4", x"aed2", x"aecf", 
    x"aecd", x"aeca", x"aec8", x"aec6", x"aec3", x"aec1", x"aebe", x"aebc", 
    x"aeb9", x"aeb7", x"aeb5", x"aeb2", x"aeb0", x"aead", x"aeab", x"aea8", 
    x"aea6", x"aea4", x"aea1", x"ae9f", x"ae9c", x"ae9a", x"ae97", x"ae95", 
    x"ae93", x"ae90", x"ae8e", x"ae8b", x"ae89", x"ae86", x"ae84", x"ae82", 
    x"ae7f", x"ae7d", x"ae7a", x"ae78", x"ae76", x"ae73", x"ae71", x"ae6e", 
    x"ae6c", x"ae69", x"ae67", x"ae65", x"ae62", x"ae60", x"ae5d", x"ae5b", 
    x"ae58", x"ae56", x"ae54", x"ae51", x"ae4f", x"ae4c", x"ae4a", x"ae48", 
    x"ae45", x"ae43", x"ae40", x"ae3e", x"ae3b", x"ae39", x"ae37", x"ae34", 
    x"ae32", x"ae2f", x"ae2d", x"ae2b", x"ae28", x"ae26", x"ae23", x"ae21", 
    x"ae1e", x"ae1c", x"ae1a", x"ae17", x"ae15", x"ae12", x"ae10", x"ae0e", 
    x"ae0b", x"ae09", x"ae06", x"ae04", x"ae02", x"adff", x"adfd", x"adfa", 
    x"adf8", x"adf5", x"adf3", x"adf1", x"adee", x"adec", x"ade9", x"ade7", 
    x"ade5", x"ade2", x"ade0", x"addd", x"addb", x"add9", x"add6", x"add4", 
    x"add1", x"adcf", x"adcd", x"adca", x"adc8", x"adc5", x"adc3", x"adc0", 
    x"adbe", x"adbc", x"adb9", x"adb7", x"adb4", x"adb2", x"adb0", x"adad", 
    x"adab", x"ada8", x"ada6", x"ada4", x"ada1", x"ad9f", x"ad9c", x"ad9a", 
    x"ad98", x"ad95", x"ad93", x"ad90", x"ad8e", x"ad8c", x"ad89", x"ad87", 
    x"ad84", x"ad82", x"ad80", x"ad7d", x"ad7b", x"ad78", x"ad76", x"ad74", 
    x"ad71", x"ad6f", x"ad6c", x"ad6a", x"ad68", x"ad65", x"ad63", x"ad60", 
    x"ad5e", x"ad5c", x"ad59", x"ad57", x"ad54", x"ad52", x"ad50", x"ad4d", 
    x"ad4b", x"ad48", x"ad46", x"ad44", x"ad41", x"ad3f", x"ad3c", x"ad3a", 
    x"ad38", x"ad35", x"ad33", x"ad30", x"ad2e", x"ad2c", x"ad29", x"ad27", 
    x"ad24", x"ad22", x"ad20", x"ad1d", x"ad1b", x"ad18", x"ad16", x"ad14", 
    x"ad11", x"ad0f", x"ad0c", x"ad0a", x"ad08", x"ad05", x"ad03", x"ad01", 
    x"acfe", x"acfc", x"acf9", x"acf7", x"acf5", x"acf2", x"acf0", x"aced", 
    x"aceb", x"ace9", x"ace6", x"ace4", x"ace1", x"acdf", x"acdd", x"acda", 
    x"acd8", x"acd6", x"acd3", x"acd1", x"acce", x"accc", x"acca", x"acc7", 
    x"acc5", x"acc2", x"acc0", x"acbe", x"acbb", x"acb9", x"acb6", x"acb4", 
    x"acb2", x"acaf", x"acad", x"acab", x"aca8", x"aca6", x"aca3", x"aca1", 
    x"ac9f", x"ac9c", x"ac9a", x"ac97", x"ac95", x"ac93", x"ac90", x"ac8e", 
    x"ac8c", x"ac89", x"ac87", x"ac84", x"ac82", x"ac80", x"ac7d", x"ac7b", 
    x"ac79", x"ac76", x"ac74", x"ac71", x"ac6f", x"ac6d", x"ac6a", x"ac68", 
    x"ac65", x"ac63", x"ac61", x"ac5e", x"ac5c", x"ac5a", x"ac57", x"ac55", 
    x"ac52", x"ac50", x"ac4e", x"ac4b", x"ac49", x"ac47", x"ac44", x"ac42", 
    x"ac3f", x"ac3d", x"ac3b", x"ac38", x"ac36", x"ac34", x"ac31", x"ac2f", 
    x"ac2c", x"ac2a", x"ac28", x"ac25", x"ac23", x"ac21", x"ac1e", x"ac1c", 
    x"ac19", x"ac17", x"ac15", x"ac12", x"ac10", x"ac0e", x"ac0b", x"ac09", 
    x"ac06", x"ac04", x"ac02", x"abff", x"abfd", x"abfb", x"abf8", x"abf6", 
    x"abf4", x"abf1", x"abef", x"abec", x"abea", x"abe8", x"abe5", x"abe3", 
    x"abe1", x"abde", x"abdc", x"abd9", x"abd7", x"abd5", x"abd2", x"abd0", 
    x"abce", x"abcb", x"abc9", x"abc7", x"abc4", x"abc2", x"abbf", x"abbd", 
    x"abbb", x"abb8", x"abb6", x"abb4", x"abb1", x"abaf", x"abad", x"abaa", 
    x"aba8", x"aba5", x"aba3", x"aba1", x"ab9e", x"ab9c", x"ab9a", x"ab97", 
    x"ab95", x"ab93", x"ab90", x"ab8e", x"ab8b", x"ab89", x"ab87", x"ab84", 
    x"ab82", x"ab80", x"ab7d", x"ab7b", x"ab79", x"ab76", x"ab74", x"ab72", 
    x"ab6f", x"ab6d", x"ab6a", x"ab68", x"ab66", x"ab63", x"ab61", x"ab5f", 
    x"ab5c", x"ab5a", x"ab58", x"ab55", x"ab53", x"ab51", x"ab4e", x"ab4c", 
    x"ab49", x"ab47", x"ab45", x"ab42", x"ab40", x"ab3e", x"ab3b", x"ab39", 
    x"ab37", x"ab34", x"ab32", x"ab30", x"ab2d", x"ab2b", x"ab29", x"ab26", 
    x"ab24", x"ab21", x"ab1f", x"ab1d", x"ab1a", x"ab18", x"ab16", x"ab13", 
    x"ab11", x"ab0f", x"ab0c", x"ab0a", x"ab08", x"ab05", x"ab03", x"ab01", 
    x"aafe", x"aafc", x"aafa", x"aaf7", x"aaf5", x"aaf2", x"aaf0", x"aaee", 
    x"aaeb", x"aae9", x"aae7", x"aae4", x"aae2", x"aae0", x"aadd", x"aadb", 
    x"aad9", x"aad6", x"aad4", x"aad2", x"aacf", x"aacd", x"aacb", x"aac8", 
    x"aac6", x"aac4", x"aac1", x"aabf", x"aabd", x"aaba", x"aab8", x"aab5", 
    x"aab3", x"aab1", x"aaae", x"aaac", x"aaaa", x"aaa7", x"aaa5", x"aaa3", 
    x"aaa0", x"aa9e", x"aa9c", x"aa99", x"aa97", x"aa95", x"aa92", x"aa90", 
    x"aa8e", x"aa8b", x"aa89", x"aa87", x"aa84", x"aa82", x"aa80", x"aa7d", 
    x"aa7b", x"aa79", x"aa76", x"aa74", x"aa72", x"aa6f", x"aa6d", x"aa6b", 
    x"aa68", x"aa66", x"aa64", x"aa61", x"aa5f", x"aa5d", x"aa5a", x"aa58", 
    x"aa56", x"aa53", x"aa51", x"aa4f", x"aa4c", x"aa4a", x"aa48", x"aa45", 
    x"aa43", x"aa41", x"aa3e", x"aa3c", x"aa3a", x"aa37", x"aa35", x"aa33", 
    x"aa30", x"aa2e", x"aa2c", x"aa29", x"aa27", x"aa25", x"aa22", x"aa20", 
    x"aa1e", x"aa1b", x"aa19", x"aa17", x"aa14", x"aa12", x"aa10", x"aa0d", 
    x"aa0b", x"aa09", x"aa06", x"aa04", x"aa02", x"a9ff", x"a9fd", x"a9fb", 
    x"a9f8", x"a9f6", x"a9f4", x"a9f1", x"a9ef", x"a9ed", x"a9ea", x"a9e8", 
    x"a9e6", x"a9e3", x"a9e1", x"a9df", x"a9dd", x"a9da", x"a9d8", x"a9d6", 
    x"a9d3", x"a9d1", x"a9cf", x"a9cc", x"a9ca", x"a9c8", x"a9c5", x"a9c3", 
    x"a9c1", x"a9be", x"a9bc", x"a9ba", x"a9b7", x"a9b5", x"a9b3", x"a9b0", 
    x"a9ae", x"a9ac", x"a9a9", x"a9a7", x"a9a5", x"a9a2", x"a9a0", x"a99e", 
    x"a99c", x"a999", x"a997", x"a995", x"a992", x"a990", x"a98e", x"a98b", 
    x"a989", x"a987", x"a984", x"a982", x"a980", x"a97d", x"a97b", x"a979", 
    x"a976", x"a974", x"a972", x"a970", x"a96d", x"a96b", x"a969", x"a966", 
    x"a964", x"a962", x"a95f", x"a95d", x"a95b", x"a958", x"a956", x"a954", 
    x"a951", x"a94f", x"a94d", x"a94b", x"a948", x"a946", x"a944", x"a941", 
    x"a93f", x"a93d", x"a93a", x"a938", x"a936", x"a933", x"a931", x"a92f", 
    x"a92d", x"a92a", x"a928", x"a926", x"a923", x"a921", x"a91f", x"a91c", 
    x"a91a", x"a918", x"a915", x"a913", x"a911", x"a90f", x"a90c", x"a90a", 
    x"a908", x"a905", x"a903", x"a901", x"a8fe", x"a8fc", x"a8fa", x"a8f7", 
    x"a8f5", x"a8f3", x"a8f1", x"a8ee", x"a8ec", x"a8ea", x"a8e7", x"a8e5", 
    x"a8e3", x"a8e0", x"a8de", x"a8dc", x"a8da", x"a8d7", x"a8d5", x"a8d3", 
    x"a8d0", x"a8ce", x"a8cc", x"a8c9", x"a8c7", x"a8c5", x"a8c3", x"a8c0", 
    x"a8be", x"a8bc", x"a8b9", x"a8b7", x"a8b5", x"a8b2", x"a8b0", x"a8ae", 
    x"a8ac", x"a8a9", x"a8a7", x"a8a5", x"a8a2", x"a8a0", x"a89e", x"a89b", 
    x"a899", x"a897", x"a895", x"a892", x"a890", x"a88e", x"a88b", x"a889", 
    x"a887", x"a885", x"a882", x"a880", x"a87e", x"a87b", x"a879", x"a877", 
    x"a875", x"a872", x"a870", x"a86e", x"a86b", x"a869", x"a867", x"a864", 
    x"a862", x"a860", x"a85e", x"a85b", x"a859", x"a857", x"a854", x"a852", 
    x"a850", x"a84e", x"a84b", x"a849", x"a847", x"a844", x"a842", x"a840", 
    x"a83e", x"a83b", x"a839", x"a837", x"a834", x"a832", x"a830", x"a82e", 
    x"a82b", x"a829", x"a827", x"a824", x"a822", x"a820", x"a81e", x"a81b", 
    x"a819", x"a817", x"a814", x"a812", x"a810", x"a80e", x"a80b", x"a809", 
    x"a807", x"a804", x"a802", x"a800", x"a7fe", x"a7fb", x"a7f9", x"a7f7", 
    x"a7f4", x"a7f2", x"a7f0", x"a7ee", x"a7eb", x"a7e9", x"a7e7", x"a7e5", 
    x"a7e2", x"a7e0", x"a7de", x"a7db", x"a7d9", x"a7d7", x"a7d5", x"a7d2", 
    x"a7d0", x"a7ce", x"a7cb", x"a7c9", x"a7c7", x"a7c5", x"a7c2", x"a7c0", 
    x"a7be", x"a7bc", x"a7b9", x"a7b7", x"a7b5", x"a7b2", x"a7b0", x"a7ae", 
    x"a7ac", x"a7a9", x"a7a7", x"a7a5", x"a7a3", x"a7a0", x"a79e", x"a79c", 
    x"a799", x"a797", x"a795", x"a793", x"a790", x"a78e", x"a78c", x"a78a", 
    x"a787", x"a785", x"a783", x"a780", x"a77e", x"a77c", x"a77a", x"a777", 
    x"a775", x"a773", x"a771", x"a76e", x"a76c", x"a76a", x"a768", x"a765", 
    x"a763", x"a761", x"a75e", x"a75c", x"a75a", x"a758", x"a755", x"a753", 
    x"a751", x"a74f", x"a74c", x"a74a", x"a748", x"a746", x"a743", x"a741", 
    x"a73f", x"a73c", x"a73a", x"a738", x"a736", x"a733", x"a731", x"a72f", 
    x"a72d", x"a72a", x"a728", x"a726", x"a724", x"a721", x"a71f", x"a71d", 
    x"a71b", x"a718", x"a716", x"a714", x"a712", x"a70f", x"a70d", x"a70b", 
    x"a708", x"a706", x"a704", x"a702", x"a6ff", x"a6fd", x"a6fb", x"a6f9", 
    x"a6f6", x"a6f4", x"a6f2", x"a6f0", x"a6ed", x"a6eb", x"a6e9", x"a6e7", 
    x"a6e4", x"a6e2", x"a6e0", x"a6de", x"a6db", x"a6d9", x"a6d7", x"a6d5", 
    x"a6d2", x"a6d0", x"a6ce", x"a6cc", x"a6c9", x"a6c7", x"a6c5", x"a6c3", 
    x"a6c0", x"a6be", x"a6bc", x"a6ba", x"a6b7", x"a6b5", x"a6b3", x"a6b1", 
    x"a6ae", x"a6ac", x"a6aa", x"a6a8", x"a6a5", x"a6a3", x"a6a1", x"a69f", 
    x"a69c", x"a69a", x"a698", x"a696", x"a693", x"a691", x"a68f", x"a68d", 
    x"a68a", x"a688", x"a686", x"a684", x"a681", x"a67f", x"a67d", x"a67b", 
    x"a678", x"a676", x"a674", x"a672", x"a66f", x"a66d", x"a66b", x"a669", 
    x"a666", x"a664", x"a662", x"a660", x"a65d", x"a65b", x"a659", x"a657", 
    x"a654", x"a652", x"a650", x"a64e", x"a64b", x"a649", x"a647", x"a645", 
    x"a643", x"a640", x"a63e", x"a63c", x"a63a", x"a637", x"a635", x"a633", 
    x"a631", x"a62e", x"a62c", x"a62a", x"a628", x"a625", x"a623", x"a621", 
    x"a61f", x"a61c", x"a61a", x"a618", x"a616", x"a614", x"a611", x"a60f", 
    x"a60d", x"a60b", x"a608", x"a606", x"a604", x"a602", x"a5ff", x"a5fd", 
    x"a5fb", x"a5f9", x"a5f6", x"a5f4", x"a5f2", x"a5f0", x"a5ee", x"a5eb", 
    x"a5e9", x"a5e7", x"a5e5", x"a5e2", x"a5e0", x"a5de", x"a5dc", x"a5d9", 
    x"a5d7", x"a5d5", x"a5d3", x"a5d1", x"a5ce", x"a5cc", x"a5ca", x"a5c8", 
    x"a5c5", x"a5c3", x"a5c1", x"a5bf", x"a5bd", x"a5ba", x"a5b8", x"a5b6", 
    x"a5b4", x"a5b1", x"a5af", x"a5ad", x"a5ab", x"a5a8", x"a5a6", x"a5a4", 
    x"a5a2", x"a5a0", x"a59d", x"a59b", x"a599", x"a597", x"a594", x"a592", 
    x"a590", x"a58e", x"a58c", x"a589", x"a587", x"a585", x"a583", x"a580", 
    x"a57e", x"a57c", x"a57a", x"a578", x"a575", x"a573", x"a571", x"a56f", 
    x"a56c", x"a56a", x"a568", x"a566", x"a564", x"a561", x"a55f", x"a55d", 
    x"a55b", x"a558", x"a556", x"a554", x"a552", x"a550", x"a54d", x"a54b", 
    x"a549", x"a547", x"a545", x"a542", x"a540", x"a53e", x"a53c", x"a539", 
    x"a537", x"a535", x"a533", x"a531", x"a52e", x"a52c", x"a52a", x"a528", 
    x"a526", x"a523", x"a521", x"a51f", x"a51d", x"a51a", x"a518", x"a516", 
    x"a514", x"a512", x"a50f", x"a50d", x"a50b", x"a509", x"a507", x"a504", 
    x"a502", x"a500", x"a4fe", x"a4fc", x"a4f9", x"a4f7", x"a4f5", x"a4f3", 
    x"a4f1", x"a4ee", x"a4ec", x"a4ea", x"a4e8", x"a4e5", x"a4e3", x"a4e1", 
    x"a4df", x"a4dd", x"a4da", x"a4d8", x"a4d6", x"a4d4", x"a4d2", x"a4cf", 
    x"a4cd", x"a4cb", x"a4c9", x"a4c7", x"a4c4", x"a4c2", x"a4c0", x"a4be", 
    x"a4bc", x"a4b9", x"a4b7", x"a4b5", x"a4b3", x"a4b1", x"a4ae", x"a4ac", 
    x"a4aa", x"a4a8", x"a4a6", x"a4a3", x"a4a1", x"a49f", x"a49d", x"a49b", 
    x"a498", x"a496", x"a494", x"a492", x"a490", x"a48d", x"a48b", x"a489", 
    x"a487", x"a485", x"a482", x"a480", x"a47e", x"a47c", x"a47a", x"a477", 
    x"a475", x"a473", x"a471", x"a46f", x"a46c", x"a46a", x"a468", x"a466", 
    x"a464", x"a461", x"a45f", x"a45d", x"a45b", x"a459", x"a456", x"a454", 
    x"a452", x"a450", x"a44e", x"a44c", x"a449", x"a447", x"a445", x"a443", 
    x"a441", x"a43e", x"a43c", x"a43a", x"a438", x"a436", x"a433", x"a431", 
    x"a42f", x"a42d", x"a42b", x"a428", x"a426", x"a424", x"a422", x"a420", 
    x"a41e", x"a41b", x"a419", x"a417", x"a415", x"a413", x"a410", x"a40e", 
    x"a40c", x"a40a", x"a408", x"a406", x"a403", x"a401", x"a3ff", x"a3fd", 
    x"a3fb", x"a3f8", x"a3f6", x"a3f4", x"a3f2", x"a3f0", x"a3ed", x"a3eb", 
    x"a3e9", x"a3e7", x"a3e5", x"a3e3", x"a3e0", x"a3de", x"a3dc", x"a3da", 
    x"a3d8", x"a3d5", x"a3d3", x"a3d1", x"a3cf", x"a3cd", x"a3cb", x"a3c8", 
    x"a3c6", x"a3c4", x"a3c2", x"a3c0", x"a3be", x"a3bb", x"a3b9", x"a3b7", 
    x"a3b5", x"a3b3", x"a3b0", x"a3ae", x"a3ac", x"a3aa", x"a3a8", x"a3a6", 
    x"a3a3", x"a3a1", x"a39f", x"a39d", x"a39b", x"a399", x"a396", x"a394", 
    x"a392", x"a390", x"a38e", x"a38c", x"a389", x"a387", x"a385", x"a383", 
    x"a381", x"a37e", x"a37c", x"a37a", x"a378", x"a376", x"a374", x"a371", 
    x"a36f", x"a36d", x"a36b", x"a369", x"a367", x"a364", x"a362", x"a360", 
    x"a35e", x"a35c", x"a35a", x"a357", x"a355", x"a353", x"a351", x"a34f", 
    x"a34d", x"a34a", x"a348", x"a346", x"a344", x"a342", x"a340", x"a33d", 
    x"a33b", x"a339", x"a337", x"a335", x"a333", x"a330", x"a32e", x"a32c", 
    x"a32a", x"a328", x"a326", x"a323", x"a321", x"a31f", x"a31d", x"a31b", 
    x"a319", x"a317", x"a314", x"a312", x"a310", x"a30e", x"a30c", x"a30a", 
    x"a307", x"a305", x"a303", x"a301", x"a2ff", x"a2fd", x"a2fa", x"a2f8", 
    x"a2f6", x"a2f4", x"a2f2", x"a2f0", x"a2ed", x"a2eb", x"a2e9", x"a2e7", 
    x"a2e5", x"a2e3", x"a2e1", x"a2de", x"a2dc", x"a2da", x"a2d8", x"a2d6", 
    x"a2d4", x"a2d1", x"a2cf", x"a2cd", x"a2cb", x"a2c9", x"a2c7", x"a2c5", 
    x"a2c2", x"a2c0", x"a2be", x"a2bc", x"a2ba", x"a2b8", x"a2b5", x"a2b3", 
    x"a2b1", x"a2af", x"a2ad", x"a2ab", x"a2a9", x"a2a6", x"a2a4", x"a2a2", 
    x"a2a0", x"a29e", x"a29c", x"a29a", x"a297", x"a295", x"a293", x"a291", 
    x"a28f", x"a28d", x"a28b", x"a288", x"a286", x"a284", x"a282", x"a280", 
    x"a27e", x"a27c", x"a279", x"a277", x"a275", x"a273", x"a271", x"a26f", 
    x"a26c", x"a26a", x"a268", x"a266", x"a264", x"a262", x"a260", x"a25d", 
    x"a25b", x"a259", x"a257", x"a255", x"a253", x"a251", x"a24f", x"a24c", 
    x"a24a", x"a248", x"a246", x"a244", x"a242", x"a240", x"a23d", x"a23b", 
    x"a239", x"a237", x"a235", x"a233", x"a231", x"a22e", x"a22c", x"a22a", 
    x"a228", x"a226", x"a224", x"a222", x"a21f", x"a21d", x"a21b", x"a219", 
    x"a217", x"a215", x"a213", x"a211", x"a20e", x"a20c", x"a20a", x"a208", 
    x"a206", x"a204", x"a202", x"a1ff", x"a1fd", x"a1fb", x"a1f9", x"a1f7", 
    x"a1f5", x"a1f3", x"a1f1", x"a1ee", x"a1ec", x"a1ea", x"a1e8", x"a1e6", 
    x"a1e4", x"a1e2", x"a1e0", x"a1dd", x"a1db", x"a1d9", x"a1d7", x"a1d5", 
    x"a1d3", x"a1d1", x"a1ce", x"a1cc", x"a1ca", x"a1c8", x"a1c6", x"a1c4", 
    x"a1c2", x"a1c0", x"a1bd", x"a1bb", x"a1b9", x"a1b7", x"a1b5", x"a1b3", 
    x"a1b1", x"a1af", x"a1ac", x"a1aa", x"a1a8", x"a1a6", x"a1a4", x"a1a2", 
    x"a1a0", x"a19e", x"a19c", x"a199", x"a197", x"a195", x"a193", x"a191", 
    x"a18f", x"a18d", x"a18b", x"a188", x"a186", x"a184", x"a182", x"a180", 
    x"a17e", x"a17c", x"a17a", x"a177", x"a175", x"a173", x"a171", x"a16f", 
    x"a16d", x"a16b", x"a169", x"a167", x"a164", x"a162", x"a160", x"a15e", 
    x"a15c", x"a15a", x"a158", x"a156", x"a153", x"a151", x"a14f", x"a14d", 
    x"a14b", x"a149", x"a147", x"a145", x"a143", x"a140", x"a13e", x"a13c", 
    x"a13a", x"a138", x"a136", x"a134", x"a132", x"a130", x"a12d", x"a12b", 
    x"a129", x"a127", x"a125", x"a123", x"a121", x"a11f", x"a11d", x"a11a", 
    x"a118", x"a116", x"a114", x"a112", x"a110", x"a10e", x"a10c", x"a10a", 
    x"a108", x"a105", x"a103", x"a101", x"a0ff", x"a0fd", x"a0fb", x"a0f9", 
    x"a0f7", x"a0f5", x"a0f2", x"a0f0", x"a0ee", x"a0ec", x"a0ea", x"a0e8", 
    x"a0e6", x"a0e4", x"a0e2", x"a0e0", x"a0dd", x"a0db", x"a0d9", x"a0d7", 
    x"a0d5", x"a0d3", x"a0d1", x"a0cf", x"a0cd", x"a0cb", x"a0c8", x"a0c6", 
    x"a0c4", x"a0c2", x"a0c0", x"a0be", x"a0bc", x"a0ba", x"a0b8", x"a0b6", 
    x"a0b3", x"a0b1", x"a0af", x"a0ad", x"a0ab", x"a0a9", x"a0a7", x"a0a5", 
    x"a0a3", x"a0a1", x"a09f", x"a09c", x"a09a", x"a098", x"a096", x"a094", 
    x"a092", x"a090", x"a08e", x"a08c", x"a08a", x"a087", x"a085", x"a083", 
    x"a081", x"a07f", x"a07d", x"a07b", x"a079", x"a077", x"a075", x"a073", 
    x"a070", x"a06e", x"a06c", x"a06a", x"a068", x"a066", x"a064", x"a062", 
    x"a060", x"a05e", x"a05c", x"a059", x"a057", x"a055", x"a053", x"a051", 
    x"a04f", x"a04d", x"a04b", x"a049", x"a047", x"a045", x"a043", x"a040", 
    x"a03e", x"a03c", x"a03a", x"a038", x"a036", x"a034", x"a032", x"a030", 
    x"a02e", x"a02c", x"a02a", x"a027", x"a025", x"a023", x"a021", x"a01f", 
    x"a01d", x"a01b", x"a019", x"a017", x"a015", x"a013", x"a011", x"a00e", 
    x"a00c", x"a00a", x"a008", x"a006", x"a004", x"a002", x"a000", x"9ffe", 
    x"9ffc", x"9ffa", x"9ff8", x"9ff6", x"9ff3", x"9ff1", x"9fef", x"9fed", 
    x"9feb", x"9fe9", x"9fe7", x"9fe5", x"9fe3", x"9fe1", x"9fdf", x"9fdd", 
    x"9fdb", x"9fd8", x"9fd6", x"9fd4", x"9fd2", x"9fd0", x"9fce", x"9fcc", 
    x"9fca", x"9fc8", x"9fc6", x"9fc4", x"9fc2", x"9fc0", x"9fbe", x"9fbb", 
    x"9fb9", x"9fb7", x"9fb5", x"9fb3", x"9fb1", x"9faf", x"9fad", x"9fab", 
    x"9fa9", x"9fa7", x"9fa5", x"9fa3", x"9fa1", x"9f9f", x"9f9c", x"9f9a", 
    x"9f98", x"9f96", x"9f94", x"9f92", x"9f90", x"9f8e", x"9f8c", x"9f8a", 
    x"9f88", x"9f86", x"9f84", x"9f82", x"9f80", x"9f7d", x"9f7b", x"9f79", 
    x"9f77", x"9f75", x"9f73", x"9f71", x"9f6f", x"9f6d", x"9f6b", x"9f69", 
    x"9f67", x"9f65", x"9f63", x"9f61", x"9f5f", x"9f5c", x"9f5a", x"9f58", 
    x"9f56", x"9f54", x"9f52", x"9f50", x"9f4e", x"9f4c", x"9f4a", x"9f48", 
    x"9f46", x"9f44", x"9f42", x"9f40", x"9f3e", x"9f3c", x"9f3a", x"9f37", 
    x"9f35", x"9f33", x"9f31", x"9f2f", x"9f2d", x"9f2b", x"9f29", x"9f27", 
    x"9f25", x"9f23", x"9f21", x"9f1f", x"9f1d", x"9f1b", x"9f19", x"9f17", 
    x"9f15", x"9f12", x"9f10", x"9f0e", x"9f0c", x"9f0a", x"9f08", x"9f06", 
    x"9f04", x"9f02", x"9f00", x"9efe", x"9efc", x"9efa", x"9ef8", x"9ef6", 
    x"9ef4", x"9ef2", x"9ef0", x"9eee", x"9eec", x"9ee9", x"9ee7", x"9ee5", 
    x"9ee3", x"9ee1", x"9edf", x"9edd", x"9edb", x"9ed9", x"9ed7", x"9ed5", 
    x"9ed3", x"9ed1", x"9ecf", x"9ecd", x"9ecb", x"9ec9", x"9ec7", x"9ec5", 
    x"9ec3", x"9ec1", x"9ebf", x"9ebd", x"9eba", x"9eb8", x"9eb6", x"9eb4", 
    x"9eb2", x"9eb0", x"9eae", x"9eac", x"9eaa", x"9ea8", x"9ea6", x"9ea4", 
    x"9ea2", x"9ea0", x"9e9e", x"9e9c", x"9e9a", x"9e98", x"9e96", x"9e94", 
    x"9e92", x"9e90", x"9e8e", x"9e8c", x"9e8a", x"9e87", x"9e85", x"9e83", 
    x"9e81", x"9e7f", x"9e7d", x"9e7b", x"9e79", x"9e77", x"9e75", x"9e73", 
    x"9e71", x"9e6f", x"9e6d", x"9e6b", x"9e69", x"9e67", x"9e65", x"9e63", 
    x"9e61", x"9e5f", x"9e5d", x"9e5b", x"9e59", x"9e57", x"9e55", x"9e53", 
    x"9e51", x"9e4f", x"9e4d", x"9e4b", x"9e48", x"9e46", x"9e44", x"9e42", 
    x"9e40", x"9e3e", x"9e3c", x"9e3a", x"9e38", x"9e36", x"9e34", x"9e32", 
    x"9e30", x"9e2e", x"9e2c", x"9e2a", x"9e28", x"9e26", x"9e24", x"9e22", 
    x"9e20", x"9e1e", x"9e1c", x"9e1a", x"9e18", x"9e16", x"9e14", x"9e12", 
    x"9e10", x"9e0e", x"9e0c", x"9e0a", x"9e08", x"9e06", x"9e04", x"9e02", 
    x"9e00", x"9dfe", x"9dfc", x"9dfa", x"9df8", x"9df5", x"9df3", x"9df1", 
    x"9def", x"9ded", x"9deb", x"9de9", x"9de7", x"9de5", x"9de3", x"9de1", 
    x"9ddf", x"9ddd", x"9ddb", x"9dd9", x"9dd7", x"9dd5", x"9dd3", x"9dd1", 
    x"9dcf", x"9dcd", x"9dcb", x"9dc9", x"9dc7", x"9dc5", x"9dc3", x"9dc1", 
    x"9dbf", x"9dbd", x"9dbb", x"9db9", x"9db7", x"9db5", x"9db3", x"9db1", 
    x"9daf", x"9dad", x"9dab", x"9da9", x"9da7", x"9da5", x"9da3", x"9da1", 
    x"9d9f", x"9d9d", x"9d9b", x"9d99", x"9d97", x"9d95", x"9d93", x"9d91", 
    x"9d8f", x"9d8d", x"9d8b", x"9d89", x"9d87", x"9d85", x"9d83", x"9d81", 
    x"9d7f", x"9d7d", x"9d7b", x"9d79", x"9d77", x"9d75", x"9d73", x"9d71", 
    x"9d6f", x"9d6d", x"9d6b", x"9d69", x"9d67", x"9d65", x"9d63", x"9d61", 
    x"9d5f", x"9d5d", x"9d5b", x"9d59", x"9d57", x"9d55", x"9d53", x"9d51", 
    x"9d4f", x"9d4d", x"9d4b", x"9d49", x"9d47", x"9d45", x"9d43", x"9d41", 
    x"9d3f", x"9d3d", x"9d3b", x"9d39", x"9d37", x"9d35", x"9d33", x"9d31", 
    x"9d2f", x"9d2d", x"9d2b", x"9d29", x"9d27", x"9d25", x"9d23", x"9d21", 
    x"9d1f", x"9d1d", x"9d1b", x"9d19", x"9d17", x"9d15", x"9d13", x"9d11", 
    x"9d0f", x"9d0d", x"9d0b", x"9d09", x"9d07", x"9d05", x"9d03", x"9d01", 
    x"9cff", x"9cfd", x"9cfb", x"9cf9", x"9cf7", x"9cf5", x"9cf3", x"9cf1", 
    x"9cef", x"9ced", x"9ceb", x"9ce9", x"9ce7", x"9ce5", x"9ce3", x"9ce1", 
    x"9cdf", x"9cdd", x"9cdb", x"9cd9", x"9cd7", x"9cd5", x"9cd3", x"9cd1", 
    x"9ccf", x"9ccd", x"9ccb", x"9cc9", x"9cc7", x"9cc5", x"9cc3", x"9cc1", 
    x"9cbf", x"9cbd", x"9cbb", x"9cb9", x"9cb7", x"9cb5", x"9cb3", x"9cb1", 
    x"9caf", x"9cad", x"9cab", x"9ca9", x"9ca7", x"9ca5", x"9ca3", x"9ca2", 
    x"9ca0", x"9c9e", x"9c9c", x"9c9a", x"9c98", x"9c96", x"9c94", x"9c92", 
    x"9c90", x"9c8e", x"9c8c", x"9c8a", x"9c88", x"9c86", x"9c84", x"9c82", 
    x"9c80", x"9c7e", x"9c7c", x"9c7a", x"9c78", x"9c76", x"9c74", x"9c72", 
    x"9c70", x"9c6e", x"9c6c", x"9c6a", x"9c68", x"9c66", x"9c64", x"9c62", 
    x"9c60", x"9c5e", x"9c5c", x"9c5a", x"9c58", x"9c56", x"9c54", x"9c52", 
    x"9c51", x"9c4f", x"9c4d", x"9c4b", x"9c49", x"9c47", x"9c45", x"9c43", 
    x"9c41", x"9c3f", x"9c3d", x"9c3b", x"9c39", x"9c37", x"9c35", x"9c33", 
    x"9c31", x"9c2f", x"9c2d", x"9c2b", x"9c29", x"9c27", x"9c25", x"9c23", 
    x"9c21", x"9c1f", x"9c1d", x"9c1b", x"9c19", x"9c17", x"9c16", x"9c14", 
    x"9c12", x"9c10", x"9c0e", x"9c0c", x"9c0a", x"9c08", x"9c06", x"9c04", 
    x"9c02", x"9c00", x"9bfe", x"9bfc", x"9bfa", x"9bf8", x"9bf6", x"9bf4", 
    x"9bf2", x"9bf0", x"9bee", x"9bec", x"9bea", x"9be8", x"9be6", x"9be4", 
    x"9be3", x"9be1", x"9bdf", x"9bdd", x"9bdb", x"9bd9", x"9bd7", x"9bd5", 
    x"9bd3", x"9bd1", x"9bcf", x"9bcd", x"9bcb", x"9bc9", x"9bc7", x"9bc5", 
    x"9bc3", x"9bc1", x"9bbf", x"9bbd", x"9bbb", x"9bb9", x"9bb8", x"9bb6", 
    x"9bb4", x"9bb2", x"9bb0", x"9bae", x"9bac", x"9baa", x"9ba8", x"9ba6", 
    x"9ba4", x"9ba2", x"9ba0", x"9b9e", x"9b9c", x"9b9a", x"9b98", x"9b96", 
    x"9b94", x"9b92", x"9b91", x"9b8f", x"9b8d", x"9b8b", x"9b89", x"9b87", 
    x"9b85", x"9b83", x"9b81", x"9b7f", x"9b7d", x"9b7b", x"9b79", x"9b77", 
    x"9b75", x"9b73", x"9b71", x"9b6f", x"9b6e", x"9b6c", x"9b6a", x"9b68", 
    x"9b66", x"9b64", x"9b62", x"9b60", x"9b5e", x"9b5c", x"9b5a", x"9b58", 
    x"9b56", x"9b54", x"9b52", x"9b50", x"9b4e", x"9b4d", x"9b4b", x"9b49", 
    x"9b47", x"9b45", x"9b43", x"9b41", x"9b3f", x"9b3d", x"9b3b", x"9b39", 
    x"9b37", x"9b35", x"9b33", x"9b31", x"9b2f", x"9b2e", x"9b2c", x"9b2a", 
    x"9b28", x"9b26", x"9b24", x"9b22", x"9b20", x"9b1e", x"9b1c", x"9b1a", 
    x"9b18", x"9b16", x"9b14", x"9b12", x"9b11", x"9b0f", x"9b0d", x"9b0b", 
    x"9b09", x"9b07", x"9b05", x"9b03", x"9b01", x"9aff", x"9afd", x"9afb", 
    x"9af9", x"9af7", x"9af6", x"9af4", x"9af2", x"9af0", x"9aee", x"9aec", 
    x"9aea", x"9ae8", x"9ae6", x"9ae4", x"9ae2", x"9ae0", x"9ade", x"9adc", 
    x"9adb", x"9ad9", x"9ad7", x"9ad5", x"9ad3", x"9ad1", x"9acf", x"9acd", 
    x"9acb", x"9ac9", x"9ac7", x"9ac5", x"9ac3", x"9ac2", x"9ac0", x"9abe", 
    x"9abc", x"9aba", x"9ab8", x"9ab6", x"9ab4", x"9ab2", x"9ab0", x"9aae", 
    x"9aac", x"9aaa", x"9aa9", x"9aa7", x"9aa5", x"9aa3", x"9aa1", x"9a9f", 
    x"9a9d", x"9a9b", x"9a99", x"9a97", x"9a95", x"9a93", x"9a92", x"9a90", 
    x"9a8e", x"9a8c", x"9a8a", x"9a88", x"9a86", x"9a84", x"9a82", x"9a80", 
    x"9a7e", x"9a7c", x"9a7b", x"9a79", x"9a77", x"9a75", x"9a73", x"9a71", 
    x"9a6f", x"9a6d", x"9a6b", x"9a69", x"9a67", x"9a66", x"9a64", x"9a62", 
    x"9a60", x"9a5e", x"9a5c", x"9a5a", x"9a58", x"9a56", x"9a54", x"9a52", 
    x"9a51", x"9a4f", x"9a4d", x"9a4b", x"9a49", x"9a47", x"9a45", x"9a43", 
    x"9a41", x"9a3f", x"9a3d", x"9a3c", x"9a3a", x"9a38", x"9a36", x"9a34", 
    x"9a32", x"9a30", x"9a2e", x"9a2c", x"9a2a", x"9a29", x"9a27", x"9a25", 
    x"9a23", x"9a21", x"9a1f", x"9a1d", x"9a1b", x"9a19", x"9a17", x"9a16", 
    x"9a14", x"9a12", x"9a10", x"9a0e", x"9a0c", x"9a0a", x"9a08", x"9a06", 
    x"9a04", x"9a03", x"9a01", x"99ff", x"99fd", x"99fb", x"99f9", x"99f7", 
    x"99f5", x"99f3", x"99f1", x"99f0", x"99ee", x"99ec", x"99ea", x"99e8", 
    x"99e6", x"99e4", x"99e2", x"99e0", x"99de", x"99dd", x"99db", x"99d9", 
    x"99d7", x"99d5", x"99d3", x"99d1", x"99cf", x"99cd", x"99cc", x"99ca", 
    x"99c8", x"99c6", x"99c4", x"99c2", x"99c0", x"99be", x"99bc", x"99bb", 
    x"99b9", x"99b7", x"99b5", x"99b3", x"99b1", x"99af", x"99ad", x"99ab", 
    x"99aa", x"99a8", x"99a6", x"99a4", x"99a2", x"99a0", x"999e", x"999c", 
    x"999a", x"9999", x"9997", x"9995", x"9993", x"9991", x"998f", x"998d", 
    x"998b", x"998a", x"9988", x"9986", x"9984", x"9982", x"9980", x"997e", 
    x"997c", x"997a", x"9979", x"9977", x"9975", x"9973", x"9971", x"996f", 
    x"996d", x"996b", x"996a", x"9968", x"9966", x"9964", x"9962", x"9960", 
    x"995e", x"995c", x"995b", x"9959", x"9957", x"9955", x"9953", x"9951", 
    x"994f", x"994d", x"994c", x"994a", x"9948", x"9946", x"9944", x"9942", 
    x"9940", x"993e", x"993d", x"993b", x"9939", x"9937", x"9935", x"9933", 
    x"9931", x"992f", x"992e", x"992c", x"992a", x"9928", x"9926", x"9924", 
    x"9922", x"9920", x"991f", x"991d", x"991b", x"9919", x"9917", x"9915", 
    x"9913", x"9912", x"9910", x"990e", x"990c", x"990a", x"9908", x"9906", 
    x"9904", x"9903", x"9901", x"98ff", x"98fd", x"98fb", x"98f9", x"98f7", 
    x"98f6", x"98f4", x"98f2", x"98f0", x"98ee", x"98ec", x"98ea", x"98e8", 
    x"98e7", x"98e5", x"98e3", x"98e1", x"98df", x"98dd", x"98db", x"98da", 
    x"98d8", x"98d6", x"98d4", x"98d2", x"98d0", x"98ce", x"98cd", x"98cb", 
    x"98c9", x"98c7", x"98c5", x"98c3", x"98c1", x"98c0", x"98be", x"98bc", 
    x"98ba", x"98b8", x"98b6", x"98b4", x"98b3", x"98b1", x"98af", x"98ad", 
    x"98ab", x"98a9", x"98a7", x"98a6", x"98a4", x"98a2", x"98a0", x"989e", 
    x"989c", x"989b", x"9899", x"9897", x"9895", x"9893", x"9891", x"988f", 
    x"988e", x"988c", x"988a", x"9888", x"9886", x"9884", x"9882", x"9881", 
    x"987f", x"987d", x"987b", x"9879", x"9877", x"9876", x"9874", x"9872", 
    x"9870", x"986e", x"986c", x"986a", x"9869", x"9867", x"9865", x"9863", 
    x"9861", x"985f", x"985e", x"985c", x"985a", x"9858", x"9856", x"9854", 
    x"9852", x"9851", x"984f", x"984d", x"984b", x"9849", x"9847", x"9846", 
    x"9844", x"9842", x"9840", x"983e", x"983c", x"983b", x"9839", x"9837", 
    x"9835", x"9833", x"9831", x"9830", x"982e", x"982c", x"982a", x"9828", 
    x"9826", x"9824", x"9823", x"9821", x"981f", x"981d", x"981b", x"9819", 
    x"9818", x"9816", x"9814", x"9812", x"9810", x"980e", x"980d", x"980b", 
    x"9809", x"9807", x"9805", x"9803", x"9802", x"9800", x"97fe", x"97fc", 
    x"97fa", x"97f9", x"97f7", x"97f5", x"97f3", x"97f1", x"97ef", x"97ee", 
    x"97ec", x"97ea", x"97e8", x"97e6", x"97e4", x"97e3", x"97e1", x"97df", 
    x"97dd", x"97db", x"97d9", x"97d8", x"97d6", x"97d4", x"97d2", x"97d0", 
    x"97ce", x"97cd", x"97cb", x"97c9", x"97c7", x"97c5", x"97c4", x"97c2", 
    x"97c0", x"97be", x"97bc", x"97ba", x"97b9", x"97b7", x"97b5", x"97b3", 
    x"97b1", x"97af", x"97ae", x"97ac", x"97aa", x"97a8", x"97a6", x"97a5", 
    x"97a3", x"97a1", x"979f", x"979d", x"979b", x"979a", x"9798", x"9796", 
    x"9794", x"9792", x"9791", x"978f", x"978d", x"978b", x"9789", x"9787", 
    x"9786", x"9784", x"9782", x"9780", x"977e", x"977d", x"977b", x"9779", 
    x"9777", x"9775", x"9774", x"9772", x"9770", x"976e", x"976c", x"976a", 
    x"9769", x"9767", x"9765", x"9763", x"9761", x"9760", x"975e", x"975c", 
    x"975a", x"9758", x"9757", x"9755", x"9753", x"9751", x"974f", x"974e", 
    x"974c", x"974a", x"9748", x"9746", x"9745", x"9743", x"9741", x"973f", 
    x"973d", x"973b", x"973a", x"9738", x"9736", x"9734", x"9732", x"9731", 
    x"972f", x"972d", x"972b", x"9729", x"9728", x"9726", x"9724", x"9722", 
    x"9720", x"971f", x"971d", x"971b", x"9719", x"9717", x"9716", x"9714", 
    x"9712", x"9710", x"970e", x"970d", x"970b", x"9709", x"9707", x"9705", 
    x"9704", x"9702", x"9700", x"96fe", x"96fc", x"96fb", x"96f9", x"96f7", 
    x"96f5", x"96f3", x"96f2", x"96f0", x"96ee", x"96ec", x"96eb", x"96e9", 
    x"96e7", x"96e5", x"96e3", x"96e2", x"96e0", x"96de", x"96dc", x"96da", 
    x"96d9", x"96d7", x"96d5", x"96d3", x"96d1", x"96d0", x"96ce", x"96cc", 
    x"96ca", x"96c8", x"96c7", x"96c5", x"96c3", x"96c1", x"96c0", x"96be", 
    x"96bc", x"96ba", x"96b8", x"96b7", x"96b5", x"96b3", x"96b1", x"96af", 
    x"96ae", x"96ac", x"96aa", x"96a8", x"96a7", x"96a5", x"96a3", x"96a1", 
    x"969f", x"969e", x"969c", x"969a", x"9698", x"9696", x"9695", x"9693", 
    x"9691", x"968f", x"968e", x"968c", x"968a", x"9688", x"9686", x"9685", 
    x"9683", x"9681", x"967f", x"967e", x"967c", x"967a", x"9678", x"9676", 
    x"9675", x"9673", x"9671", x"966f", x"966e", x"966c", x"966a", x"9668", 
    x"9666", x"9665", x"9663", x"9661", x"965f", x"965e", x"965c", x"965a", 
    x"9658", x"9657", x"9655", x"9653", x"9651", x"964f", x"964e", x"964c", 
    x"964a", x"9648", x"9647", x"9645", x"9643", x"9641", x"963f", x"963e", 
    x"963c", x"963a", x"9638", x"9637", x"9635", x"9633", x"9631", x"9630", 
    x"962e", x"962c", x"962a", x"9628", x"9627", x"9625", x"9623", x"9621", 
    x"9620", x"961e", x"961c", x"961a", x"9619", x"9617", x"9615", x"9613", 
    x"9612", x"9610", x"960e", x"960c", x"960a", x"9609", x"9607", x"9605", 
    x"9603", x"9602", x"9600", x"95fe", x"95fc", x"95fb", x"95f9", x"95f7", 
    x"95f5", x"95f4", x"95f2", x"95f0", x"95ee", x"95ed", x"95eb", x"95e9", 
    x"95e7", x"95e6", x"95e4", x"95e2", x"95e0", x"95df", x"95dd", x"95db", 
    x"95d9", x"95d7", x"95d6", x"95d4", x"95d2", x"95d0", x"95cf", x"95cd", 
    x"95cb", x"95c9", x"95c8", x"95c6", x"95c4", x"95c2", x"95c1", x"95bf", 
    x"95bd", x"95bb", x"95ba", x"95b8", x"95b6", x"95b4", x"95b3", x"95b1", 
    x"95af", x"95ad", x"95ac", x"95aa", x"95a8", x"95a6", x"95a5", x"95a3", 
    x"95a1", x"959f", x"959e", x"959c", x"959a", x"9598", x"9597", x"9595", 
    x"9593", x"9591", x"9590", x"958e", x"958c", x"958b", x"9589", x"9587", 
    x"9585", x"9584", x"9582", x"9580", x"957e", x"957d", x"957b", x"9579", 
    x"9577", x"9576", x"9574", x"9572", x"9570", x"956f", x"956d", x"956b", 
    x"9569", x"9568", x"9566", x"9564", x"9562", x"9561", x"955f", x"955d", 
    x"955c", x"955a", x"9558", x"9556", x"9555", x"9553", x"9551", x"954f", 
    x"954e", x"954c", x"954a", x"9548", x"9547", x"9545", x"9543", x"9541", 
    x"9540", x"953e", x"953c", x"953b", x"9539", x"9537", x"9535", x"9534", 
    x"9532", x"9530", x"952e", x"952d", x"952b", x"9529", x"9528", x"9526", 
    x"9524", x"9522", x"9521", x"951f", x"951d", x"951b", x"951a", x"9518", 
    x"9516", x"9514", x"9513", x"9511", x"950f", x"950e", x"950c", x"950a", 
    x"9508", x"9507", x"9505", x"9503", x"9502", x"9500", x"94fe", x"94fc", 
    x"94fb", x"94f9", x"94f7", x"94f5", x"94f4", x"94f2", x"94f0", x"94ef", 
    x"94ed", x"94eb", x"94e9", x"94e8", x"94e6", x"94e4", x"94e3", x"94e1", 
    x"94df", x"94dd", x"94dc", x"94da", x"94d8", x"94d6", x"94d5", x"94d3", 
    x"94d1", x"94d0", x"94ce", x"94cc", x"94ca", x"94c9", x"94c7", x"94c5", 
    x"94c4", x"94c2", x"94c0", x"94be", x"94bd", x"94bb", x"94b9", x"94b8", 
    x"94b6", x"94b4", x"94b2", x"94b1", x"94af", x"94ad", x"94ac", x"94aa", 
    x"94a8", x"94a6", x"94a5", x"94a3", x"94a1", x"94a0", x"949e", x"949c", 
    x"949b", x"9499", x"9497", x"9495", x"9494", x"9492", x"9490", x"948f", 
    x"948d", x"948b", x"9489", x"9488", x"9486", x"9484", x"9483", x"9481", 
    x"947f", x"947d", x"947c", x"947a", x"9478", x"9477", x"9475", x"9473", 
    x"9472", x"9470", x"946e", x"946c", x"946b", x"9469", x"9467", x"9466", 
    x"9464", x"9462", x"9461", x"945f", x"945d", x"945b", x"945a", x"9458", 
    x"9456", x"9455", x"9453", x"9451", x"9450", x"944e", x"944c", x"944a", 
    x"9449", x"9447", x"9445", x"9444", x"9442", x"9440", x"943f", x"943d", 
    x"943b", x"943a", x"9438", x"9436", x"9434", x"9433", x"9431", x"942f", 
    x"942e", x"942c", x"942a", x"9429", x"9427", x"9425", x"9423", x"9422", 
    x"9420", x"941e", x"941d", x"941b", x"9419", x"9418", x"9416", x"9414", 
    x"9413", x"9411", x"940f", x"940e", x"940c", x"940a", x"9408", x"9407", 
    x"9405", x"9403", x"9402", x"9400", x"93fe", x"93fd", x"93fb", x"93f9", 
    x"93f8", x"93f6", x"93f4", x"93f3", x"93f1", x"93ef", x"93ee", x"93ec", 
    x"93ea", x"93e8", x"93e7", x"93e5", x"93e3", x"93e2", x"93e0", x"93de", 
    x"93dd", x"93db", x"93d9", x"93d8", x"93d6", x"93d4", x"93d3", x"93d1", 
    x"93cf", x"93ce", x"93cc", x"93ca", x"93c9", x"93c7", x"93c5", x"93c4", 
    x"93c2", x"93c0", x"93be", x"93bd", x"93bb", x"93b9", x"93b8", x"93b6", 
    x"93b4", x"93b3", x"93b1", x"93af", x"93ae", x"93ac", x"93aa", x"93a9", 
    x"93a7", x"93a5", x"93a4", x"93a2", x"93a0", x"939f", x"939d", x"939b", 
    x"939a", x"9398", x"9396", x"9395", x"9393", x"9391", x"9390", x"938e", 
    x"938c", x"938b", x"9389", x"9387", x"9386", x"9384", x"9382", x"9381", 
    x"937f", x"937d", x"937c", x"937a", x"9378", x"9377", x"9375", x"9373", 
    x"9372", x"9370", x"936e", x"936d", x"936b", x"9369", x"9368", x"9366", 
    x"9364", x"9363", x"9361", x"935f", x"935e", x"935c", x"935a", x"9359", 
    x"9357", x"9355", x"9354", x"9352", x"9350", x"934f", x"934d", x"934b", 
    x"934a", x"9348", x"9346", x"9345", x"9343", x"9341", x"9340", x"933e", 
    x"933d", x"933b", x"9339", x"9338", x"9336", x"9334", x"9333", x"9331", 
    x"932f", x"932e", x"932c", x"932a", x"9329", x"9327", x"9325", x"9324", 
    x"9322", x"9320", x"931f", x"931d", x"931b", x"931a", x"9318", x"9316", 
    x"9315", x"9313", x"9312", x"9310", x"930e", x"930d", x"930b", x"9309", 
    x"9308", x"9306", x"9304", x"9303", x"9301", x"92ff", x"92fe", x"92fc", 
    x"92fa", x"92f9", x"92f7", x"92f6", x"92f4", x"92f2", x"92f1", x"92ef", 
    x"92ed", x"92ec", x"92ea", x"92e8", x"92e7", x"92e5", x"92e3", x"92e2", 
    x"92e0", x"92df", x"92dd", x"92db", x"92da", x"92d8", x"92d6", x"92d5", 
    x"92d3", x"92d1", x"92d0", x"92ce", x"92cc", x"92cb", x"92c9", x"92c8", 
    x"92c6", x"92c4", x"92c3", x"92c1", x"92bf", x"92be", x"92bc", x"92ba", 
    x"92b9", x"92b7", x"92b6", x"92b4", x"92b2", x"92b1", x"92af", x"92ad", 
    x"92ac", x"92aa", x"92a8", x"92a7", x"92a5", x"92a4", x"92a2", x"92a0", 
    x"929f", x"929d", x"929b", x"929a", x"9298", x"9297", x"9295", x"9293", 
    x"9292", x"9290", x"928e", x"928d", x"928b", x"928a", x"9288", x"9286", 
    x"9285", x"9283", x"9281", x"9280", x"927e", x"927c", x"927b", x"9279", 
    x"9278", x"9276", x"9274", x"9273", x"9271", x"926f", x"926e", x"926c", 
    x"926b", x"9269", x"9267", x"9266", x"9264", x"9263", x"9261", x"925f", 
    x"925e", x"925c", x"925a", x"9259", x"9257", x"9256", x"9254", x"9252", 
    x"9251", x"924f", x"924d", x"924c", x"924a", x"9249", x"9247", x"9245", 
    x"9244", x"9242", x"9241", x"923f", x"923d", x"923c", x"923a", x"9238", 
    x"9237", x"9235", x"9234", x"9232", x"9230", x"922f", x"922d", x"922c", 
    x"922a", x"9228", x"9227", x"9225", x"9223", x"9222", x"9220", x"921f", 
    x"921d", x"921b", x"921a", x"9218", x"9217", x"9215", x"9213", x"9212", 
    x"9210", x"920f", x"920d", x"920b", x"920a", x"9208", x"9206", x"9205", 
    x"9203", x"9202", x"9200", x"91fe", x"91fd", x"91fb", x"91fa", x"91f8", 
    x"91f6", x"91f5", x"91f3", x"91f2", x"91f0", x"91ee", x"91ed", x"91eb", 
    x"91ea", x"91e8", x"91e6", x"91e5", x"91e3", x"91e2", x"91e0", x"91de", 
    x"91dd", x"91db", x"91da", x"91d8", x"91d6", x"91d5", x"91d3", x"91d2", 
    x"91d0", x"91ce", x"91cd", x"91cb", x"91ca", x"91c8", x"91c6", x"91c5", 
    x"91c3", x"91c2", x"91c0", x"91be", x"91bd", x"91bb", x"91ba", x"91b8", 
    x"91b6", x"91b5", x"91b3", x"91b2", x"91b0", x"91ae", x"91ad", x"91ab", 
    x"91aa", x"91a8", x"91a7", x"91a5", x"91a3", x"91a2", x"91a0", x"919f", 
    x"919d", x"919b", x"919a", x"9198", x"9197", x"9195", x"9193", x"9192", 
    x"9190", x"918f", x"918d", x"918b", x"918a", x"9188", x"9187", x"9185", 
    x"9184", x"9182", x"9180", x"917f", x"917d", x"917c", x"917a", x"9178", 
    x"9177", x"9175", x"9174", x"9172", x"9171", x"916f", x"916d", x"916c", 
    x"916a", x"9169", x"9167", x"9165", x"9164", x"9162", x"9161", x"915f", 
    x"915e", x"915c", x"915a", x"9159", x"9157", x"9156", x"9154", x"9153", 
    x"9151", x"914f", x"914e", x"914c", x"914b", x"9149", x"9147", x"9146", 
    x"9144", x"9143", x"9141", x"9140", x"913e", x"913c", x"913b", x"9139", 
    x"9138", x"9136", x"9135", x"9133", x"9131", x"9130", x"912e", x"912d", 
    x"912b", x"912a", x"9128", x"9126", x"9125", x"9123", x"9122", x"9120", 
    x"911f", x"911d", x"911b", x"911a", x"9118", x"9117", x"9115", x"9114", 
    x"9112", x"9110", x"910f", x"910d", x"910c", x"910a", x"9109", x"9107", 
    x"9105", x"9104", x"9102", x"9101", x"90ff", x"90fe", x"90fc", x"90fb", 
    x"90f9", x"90f7", x"90f6", x"90f4", x"90f3", x"90f1", x"90f0", x"90ee", 
    x"90ec", x"90eb", x"90e9", x"90e8", x"90e6", x"90e5", x"90e3", x"90e2", 
    x"90e0", x"90de", x"90dd", x"90db", x"90da", x"90d8", x"90d7", x"90d5", 
    x"90d4", x"90d2", x"90d0", x"90cf", x"90cd", x"90cc", x"90ca", x"90c9", 
    x"90c7", x"90c6", x"90c4", x"90c2", x"90c1", x"90bf", x"90be", x"90bc", 
    x"90bb", x"90b9", x"90b8", x"90b6", x"90b4", x"90b3", x"90b1", x"90b0", 
    x"90ae", x"90ad", x"90ab", x"90aa", x"90a8", x"90a7", x"90a5", x"90a3", 
    x"90a2", x"90a0", x"909f", x"909d", x"909c", x"909a", x"9099", x"9097", 
    x"9095", x"9094", x"9092", x"9091", x"908f", x"908e", x"908c", x"908b", 
    x"9089", x"9088", x"9086", x"9084", x"9083", x"9081", x"9080", x"907e", 
    x"907d", x"907b", x"907a", x"9078", x"9077", x"9075", x"9074", x"9072", 
    x"9070", x"906f", x"906d", x"906c", x"906a", x"9069", x"9067", x"9066", 
    x"9064", x"9063", x"9061", x"9060", x"905e", x"905c", x"905b", x"9059", 
    x"9058", x"9056", x"9055", x"9053", x"9052", x"9050", x"904f", x"904d", 
    x"904c", x"904a", x"9048", x"9047", x"9045", x"9044", x"9042", x"9041", 
    x"903f", x"903e", x"903c", x"903b", x"9039", x"9038", x"9036", x"9035", 
    x"9033", x"9032", x"9030", x"902e", x"902d", x"902b", x"902a", x"9028", 
    x"9027", x"9025", x"9024", x"9022", x"9021", x"901f", x"901e", x"901c", 
    x"901b", x"9019", x"9018", x"9016", x"9015", x"9013", x"9011", x"9010", 
    x"900e", x"900d", x"900b", x"900a", x"9008", x"9007", x"9005", x"9004", 
    x"9002", x"9001", x"8fff", x"8ffe", x"8ffc", x"8ffb", x"8ff9", x"8ff8", 
    x"8ff6", x"8ff5", x"8ff3", x"8ff2", x"8ff0", x"8fee", x"8fed", x"8feb", 
    x"8fea", x"8fe8", x"8fe7", x"8fe5", x"8fe4", x"8fe2", x"8fe1", x"8fdf", 
    x"8fde", x"8fdc", x"8fdb", x"8fd9", x"8fd8", x"8fd6", x"8fd5", x"8fd3", 
    x"8fd2", x"8fd0", x"8fcf", x"8fcd", x"8fcc", x"8fca", x"8fc9", x"8fc7", 
    x"8fc6", x"8fc4", x"8fc3", x"8fc1", x"8fc0", x"8fbe", x"8fbd", x"8fbb", 
    x"8fba", x"8fb8", x"8fb7", x"8fb5", x"8fb4", x"8fb2", x"8fb0", x"8faf", 
    x"8fad", x"8fac", x"8faa", x"8fa9", x"8fa7", x"8fa6", x"8fa4", x"8fa3", 
    x"8fa1", x"8fa0", x"8f9e", x"8f9d", x"8f9b", x"8f9a", x"8f98", x"8f97", 
    x"8f95", x"8f94", x"8f92", x"8f91", x"8f8f", x"8f8e", x"8f8c", x"8f8b", 
    x"8f89", x"8f88", x"8f86", x"8f85", x"8f83", x"8f82", x"8f80", x"8f7f", 
    x"8f7d", x"8f7c", x"8f7a", x"8f79", x"8f77", x"8f76", x"8f74", x"8f73", 
    x"8f71", x"8f70", x"8f6e", x"8f6d", x"8f6b", x"8f6a", x"8f68", x"8f67", 
    x"8f65", x"8f64", x"8f62", x"8f61", x"8f60", x"8f5e", x"8f5d", x"8f5b", 
    x"8f5a", x"8f58", x"8f57", x"8f55", x"8f54", x"8f52", x"8f51", x"8f4f", 
    x"8f4e", x"8f4c", x"8f4b", x"8f49", x"8f48", x"8f46", x"8f45", x"8f43", 
    x"8f42", x"8f40", x"8f3f", x"8f3d", x"8f3c", x"8f3a", x"8f39", x"8f37", 
    x"8f36", x"8f34", x"8f33", x"8f31", x"8f30", x"8f2e", x"8f2d", x"8f2b", 
    x"8f2a", x"8f28", x"8f27", x"8f25", x"8f24", x"8f23", x"8f21", x"8f20", 
    x"8f1e", x"8f1d", x"8f1b", x"8f1a", x"8f18", x"8f17", x"8f15", x"8f14", 
    x"8f12", x"8f11", x"8f0f", x"8f0e", x"8f0c", x"8f0b", x"8f09", x"8f08", 
    x"8f06", x"8f05", x"8f03", x"8f02", x"8f01", x"8eff", x"8efe", x"8efc", 
    x"8efb", x"8ef9", x"8ef8", x"8ef6", x"8ef5", x"8ef3", x"8ef2", x"8ef0", 
    x"8eef", x"8eed", x"8eec", x"8eea", x"8ee9", x"8ee7", x"8ee6", x"8ee5", 
    x"8ee3", x"8ee2", x"8ee0", x"8edf", x"8edd", x"8edc", x"8eda", x"8ed9", 
    x"8ed7", x"8ed6", x"8ed4", x"8ed3", x"8ed1", x"8ed0", x"8ecf", x"8ecd", 
    x"8ecc", x"8eca", x"8ec9", x"8ec7", x"8ec6", x"8ec4", x"8ec3", x"8ec1", 
    x"8ec0", x"8ebe", x"8ebd", x"8ebb", x"8eba", x"8eb9", x"8eb7", x"8eb6", 
    x"8eb4", x"8eb3", x"8eb1", x"8eb0", x"8eae", x"8ead", x"8eab", x"8eaa", 
    x"8ea8", x"8ea7", x"8ea6", x"8ea4", x"8ea3", x"8ea1", x"8ea0", x"8e9e", 
    x"8e9d", x"8e9b", x"8e9a", x"8e98", x"8e97", x"8e96", x"8e94", x"8e93", 
    x"8e91", x"8e90", x"8e8e", x"8e8d", x"8e8b", x"8e8a", x"8e88", x"8e87", 
    x"8e86", x"8e84", x"8e83", x"8e81", x"8e80", x"8e7e", x"8e7d", x"8e7b", 
    x"8e7a", x"8e78", x"8e77", x"8e76", x"8e74", x"8e73", x"8e71", x"8e70", 
    x"8e6e", x"8e6d", x"8e6b", x"8e6a", x"8e69", x"8e67", x"8e66", x"8e64", 
    x"8e63", x"8e61", x"8e60", x"8e5e", x"8e5d", x"8e5b", x"8e5a", x"8e59", 
    x"8e57", x"8e56", x"8e54", x"8e53", x"8e51", x"8e50", x"8e4e", x"8e4d", 
    x"8e4c", x"8e4a", x"8e49", x"8e47", x"8e46", x"8e44", x"8e43", x"8e42", 
    x"8e40", x"8e3f", x"8e3d", x"8e3c", x"8e3a", x"8e39", x"8e37", x"8e36", 
    x"8e35", x"8e33", x"8e32", x"8e30", x"8e2f", x"8e2d", x"8e2c", x"8e2a", 
    x"8e29", x"8e28", x"8e26", x"8e25", x"8e23", x"8e22", x"8e20", x"8e1f", 
    x"8e1e", x"8e1c", x"8e1b", x"8e19", x"8e18", x"8e16", x"8e15", x"8e14", 
    x"8e12", x"8e11", x"8e0f", x"8e0e", x"8e0c", x"8e0b", x"8e0a", x"8e08", 
    x"8e07", x"8e05", x"8e04", x"8e02", x"8e01", x"8e00", x"8dfe", x"8dfd", 
    x"8dfb", x"8dfa", x"8df8", x"8df7", x"8df6", x"8df4", x"8df3", x"8df1", 
    x"8df0", x"8dee", x"8ded", x"8dec", x"8dea", x"8de9", x"8de7", x"8de6", 
    x"8de4", x"8de3", x"8de2", x"8de0", x"8ddf", x"8ddd", x"8ddc", x"8dda", 
    x"8dd9", x"8dd8", x"8dd6", x"8dd5", x"8dd3", x"8dd2", x"8dd1", x"8dcf", 
    x"8dce", x"8dcc", x"8dcb", x"8dc9", x"8dc8", x"8dc7", x"8dc5", x"8dc4", 
    x"8dc2", x"8dc1", x"8dc0", x"8dbe", x"8dbd", x"8dbb", x"8dba", x"8db8", 
    x"8db7", x"8db6", x"8db4", x"8db3", x"8db1", x"8db0", x"8daf", x"8dad", 
    x"8dac", x"8daa", x"8da9", x"8da7", x"8da6", x"8da5", x"8da3", x"8da2", 
    x"8da0", x"8d9f", x"8d9e", x"8d9c", x"8d9b", x"8d99", x"8d98", x"8d97", 
    x"8d95", x"8d94", x"8d92", x"8d91", x"8d90", x"8d8e", x"8d8d", x"8d8b", 
    x"8d8a", x"8d88", x"8d87", x"8d86", x"8d84", x"8d83", x"8d81", x"8d80", 
    x"8d7f", x"8d7d", x"8d7c", x"8d7a", x"8d79", x"8d78", x"8d76", x"8d75", 
    x"8d73", x"8d72", x"8d71", x"8d6f", x"8d6e", x"8d6c", x"8d6b", x"8d6a", 
    x"8d68", x"8d67", x"8d65", x"8d64", x"8d63", x"8d61", x"8d60", x"8d5e", 
    x"8d5d", x"8d5c", x"8d5a", x"8d59", x"8d57", x"8d56", x"8d55", x"8d53", 
    x"8d52", x"8d50", x"8d4f", x"8d4e", x"8d4c", x"8d4b", x"8d4a", x"8d48", 
    x"8d47", x"8d45", x"8d44", x"8d43", x"8d41", x"8d40", x"8d3e", x"8d3d", 
    x"8d3c", x"8d3a", x"8d39", x"8d37", x"8d36", x"8d35", x"8d33", x"8d32", 
    x"8d30", x"8d2f", x"8d2e", x"8d2c", x"8d2b", x"8d2a", x"8d28", x"8d27", 
    x"8d25", x"8d24", x"8d23", x"8d21", x"8d20", x"8d1e", x"8d1d", x"8d1c", 
    x"8d1a", x"8d19", x"8d18", x"8d16", x"8d15", x"8d13", x"8d12", x"8d11", 
    x"8d0f", x"8d0e", x"8d0c", x"8d0b", x"8d0a", x"8d08", x"8d07", x"8d06", 
    x"8d04", x"8d03", x"8d01", x"8d00", x"8cff", x"8cfd", x"8cfc", x"8cfb", 
    x"8cf9", x"8cf8", x"8cf6", x"8cf5", x"8cf4", x"8cf2", x"8cf1", x"8cef", 
    x"8cee", x"8ced", x"8ceb", x"8cea", x"8ce9", x"8ce7", x"8ce6", x"8ce4", 
    x"8ce3", x"8ce2", x"8ce0", x"8cdf", x"8cde", x"8cdc", x"8cdb", x"8cda", 
    x"8cd8", x"8cd7", x"8cd5", x"8cd4", x"8cd3", x"8cd1", x"8cd0", x"8ccf", 
    x"8ccd", x"8ccc", x"8cca", x"8cc9", x"8cc8", x"8cc6", x"8cc5", x"8cc4", 
    x"8cc2", x"8cc1", x"8cc0", x"8cbe", x"8cbd", x"8cbb", x"8cba", x"8cb9", 
    x"8cb7", x"8cb6", x"8cb5", x"8cb3", x"8cb2", x"8cb0", x"8caf", x"8cae", 
    x"8cac", x"8cab", x"8caa", x"8ca8", x"8ca7", x"8ca6", x"8ca4", x"8ca3", 
    x"8ca2", x"8ca0", x"8c9f", x"8c9d", x"8c9c", x"8c9b", x"8c99", x"8c98", 
    x"8c97", x"8c95", x"8c94", x"8c93", x"8c91", x"8c90", x"8c8e", x"8c8d", 
    x"8c8c", x"8c8a", x"8c89", x"8c88", x"8c86", x"8c85", x"8c84", x"8c82", 
    x"8c81", x"8c80", x"8c7e", x"8c7d", x"8c7c", x"8c7a", x"8c79", x"8c77", 
    x"8c76", x"8c75", x"8c73", x"8c72", x"8c71", x"8c6f", x"8c6e", x"8c6d", 
    x"8c6b", x"8c6a", x"8c69", x"8c67", x"8c66", x"8c65", x"8c63", x"8c62", 
    x"8c61", x"8c5f", x"8c5e", x"8c5c", x"8c5b", x"8c5a", x"8c58", x"8c57", 
    x"8c56", x"8c54", x"8c53", x"8c52", x"8c50", x"8c4f", x"8c4e", x"8c4c", 
    x"8c4b", x"8c4a", x"8c48", x"8c47", x"8c46", x"8c44", x"8c43", x"8c42", 
    x"8c40", x"8c3f", x"8c3e", x"8c3c", x"8c3b", x"8c3a", x"8c38", x"8c37", 
    x"8c36", x"8c34", x"8c33", x"8c32", x"8c30", x"8c2f", x"8c2d", x"8c2c", 
    x"8c2b", x"8c29", x"8c28", x"8c27", x"8c25", x"8c24", x"8c23", x"8c21", 
    x"8c20", x"8c1f", x"8c1d", x"8c1c", x"8c1b", x"8c19", x"8c18", x"8c17", 
    x"8c15", x"8c14", x"8c13", x"8c11", x"8c10", x"8c0f", x"8c0d", x"8c0c", 
    x"8c0b", x"8c09", x"8c08", x"8c07", x"8c06", x"8c04", x"8c03", x"8c02", 
    x"8c00", x"8bff", x"8bfe", x"8bfc", x"8bfb", x"8bfa", x"8bf8", x"8bf7", 
    x"8bf6", x"8bf4", x"8bf3", x"8bf2", x"8bf0", x"8bef", x"8bee", x"8bec", 
    x"8beb", x"8bea", x"8be8", x"8be7", x"8be6", x"8be4", x"8be3", x"8be2", 
    x"8be0", x"8bdf", x"8bde", x"8bdc", x"8bdb", x"8bda", x"8bd8", x"8bd7", 
    x"8bd6", x"8bd5", x"8bd3", x"8bd2", x"8bd1", x"8bcf", x"8bce", x"8bcd", 
    x"8bcb", x"8bca", x"8bc9", x"8bc7", x"8bc6", x"8bc5", x"8bc3", x"8bc2", 
    x"8bc1", x"8bbf", x"8bbe", x"8bbd", x"8bbc", x"8bba", x"8bb9", x"8bb8", 
    x"8bb6", x"8bb5", x"8bb4", x"8bb2", x"8bb1", x"8bb0", x"8bae", x"8bad", 
    x"8bac", x"8baa", x"8ba9", x"8ba8", x"8ba7", x"8ba5", x"8ba4", x"8ba3", 
    x"8ba1", x"8ba0", x"8b9f", x"8b9d", x"8b9c", x"8b9b", x"8b99", x"8b98", 
    x"8b97", x"8b96", x"8b94", x"8b93", x"8b92", x"8b90", x"8b8f", x"8b8e", 
    x"8b8c", x"8b8b", x"8b8a", x"8b88", x"8b87", x"8b86", x"8b85", x"8b83", 
    x"8b82", x"8b81", x"8b7f", x"8b7e", x"8b7d", x"8b7b", x"8b7a", x"8b79", 
    x"8b78", x"8b76", x"8b75", x"8b74", x"8b72", x"8b71", x"8b70", x"8b6e", 
    x"8b6d", x"8b6c", x"8b6b", x"8b69", x"8b68", x"8b67", x"8b65", x"8b64", 
    x"8b63", x"8b62", x"8b60", x"8b5f", x"8b5e", x"8b5c", x"8b5b", x"8b5a", 
    x"8b58", x"8b57", x"8b56", x"8b55", x"8b53", x"8b52", x"8b51", x"8b4f", 
    x"8b4e", x"8b4d", x"8b4c", x"8b4a", x"8b49", x"8b48", x"8b46", x"8b45", 
    x"8b44", x"8b43", x"8b41", x"8b40", x"8b3f", x"8b3d", x"8b3c", x"8b3b", 
    x"8b3a", x"8b38", x"8b37", x"8b36", x"8b34", x"8b33", x"8b32", x"8b31", 
    x"8b2f", x"8b2e", x"8b2d", x"8b2b", x"8b2a", x"8b29", x"8b28", x"8b26", 
    x"8b25", x"8b24", x"8b22", x"8b21", x"8b20", x"8b1f", x"8b1d", x"8b1c", 
    x"8b1b", x"8b19", x"8b18", x"8b17", x"8b16", x"8b14", x"8b13", x"8b12", 
    x"8b10", x"8b0f", x"8b0e", x"8b0d", x"8b0b", x"8b0a", x"8b09", x"8b08", 
    x"8b06", x"8b05", x"8b04", x"8b02", x"8b01", x"8b00", x"8aff", x"8afd", 
    x"8afc", x"8afb", x"8afa", x"8af8", x"8af7", x"8af6", x"8af4", x"8af3", 
    x"8af2", x"8af1", x"8aef", x"8aee", x"8aed", x"8aec", x"8aea", x"8ae9", 
    x"8ae8", x"8ae6", x"8ae5", x"8ae4", x"8ae3", x"8ae1", x"8ae0", x"8adf", 
    x"8ade", x"8adc", x"8adb", x"8ada", x"8ad9", x"8ad7", x"8ad6", x"8ad5", 
    x"8ad3", x"8ad2", x"8ad1", x"8ad0", x"8ace", x"8acd", x"8acc", x"8acb", 
    x"8ac9", x"8ac8", x"8ac7", x"8ac6", x"8ac4", x"8ac3", x"8ac2", x"8ac1", 
    x"8abf", x"8abe", x"8abd", x"8abc", x"8aba", x"8ab9", x"8ab8", x"8ab6", 
    x"8ab5", x"8ab4", x"8ab3", x"8ab1", x"8ab0", x"8aaf", x"8aae", x"8aac", 
    x"8aab", x"8aaa", x"8aa9", x"8aa7", x"8aa6", x"8aa5", x"8aa4", x"8aa2", 
    x"8aa1", x"8aa0", x"8a9f", x"8a9d", x"8a9c", x"8a9b", x"8a9a", x"8a98", 
    x"8a97", x"8a96", x"8a95", x"8a93", x"8a92", x"8a91", x"8a90", x"8a8e", 
    x"8a8d", x"8a8c", x"8a8b", x"8a89", x"8a88", x"8a87", x"8a86", x"8a84", 
    x"8a83", x"8a82", x"8a81", x"8a7f", x"8a7e", x"8a7d", x"8a7c", x"8a7a", 
    x"8a79", x"8a78", x"8a77", x"8a75", x"8a74", x"8a73", x"8a72", x"8a70", 
    x"8a6f", x"8a6e", x"8a6d", x"8a6c", x"8a6a", x"8a69", x"8a68", x"8a67", 
    x"8a65", x"8a64", x"8a63", x"8a62", x"8a60", x"8a5f", x"8a5e", x"8a5d", 
    x"8a5b", x"8a5a", x"8a59", x"8a58", x"8a56", x"8a55", x"8a54", x"8a53", 
    x"8a52", x"8a50", x"8a4f", x"8a4e", x"8a4d", x"8a4b", x"8a4a", x"8a49", 
    x"8a48", x"8a46", x"8a45", x"8a44", x"8a43", x"8a41", x"8a40", x"8a3f", 
    x"8a3e", x"8a3d", x"8a3b", x"8a3a", x"8a39", x"8a38", x"8a36", x"8a35", 
    x"8a34", x"8a33", x"8a31", x"8a30", x"8a2f", x"8a2e", x"8a2d", x"8a2b", 
    x"8a2a", x"8a29", x"8a28", x"8a26", x"8a25", x"8a24", x"8a23", x"8a22", 
    x"8a20", x"8a1f", x"8a1e", x"8a1d", x"8a1b", x"8a1a", x"8a19", x"8a18", 
    x"8a17", x"8a15", x"8a14", x"8a13", x"8a12", x"8a10", x"8a0f", x"8a0e", 
    x"8a0d", x"8a0c", x"8a0a", x"8a09", x"8a08", x"8a07", x"8a05", x"8a04", 
    x"8a03", x"8a02", x"8a01", x"89ff", x"89fe", x"89fd", x"89fc", x"89fa", 
    x"89f9", x"89f8", x"89f7", x"89f6", x"89f4", x"89f3", x"89f2", x"89f1", 
    x"89f0", x"89ee", x"89ed", x"89ec", x"89eb", x"89e9", x"89e8", x"89e7", 
    x"89e6", x"89e5", x"89e3", x"89e2", x"89e1", x"89e0", x"89df", x"89dd", 
    x"89dc", x"89db", x"89da", x"89d9", x"89d7", x"89d6", x"89d5", x"89d4", 
    x"89d3", x"89d1", x"89d0", x"89cf", x"89ce", x"89cc", x"89cb", x"89ca", 
    x"89c9", x"89c8", x"89c6", x"89c5", x"89c4", x"89c3", x"89c2", x"89c0", 
    x"89bf", x"89be", x"89bd", x"89bc", x"89ba", x"89b9", x"89b8", x"89b7", 
    x"89b6", x"89b4", x"89b3", x"89b2", x"89b1", x"89b0", x"89ae", x"89ad", 
    x"89ac", x"89ab", x"89aa", x"89a8", x"89a7", x"89a6", x"89a5", x"89a4", 
    x"89a2", x"89a1", x"89a0", x"899f", x"899e", x"899c", x"899b", x"899a", 
    x"8999", x"8998", x"8997", x"8995", x"8994", x"8993", x"8992", x"8991", 
    x"898f", x"898e", x"898d", x"898c", x"898b", x"8989", x"8988", x"8987", 
    x"8986", x"8985", x"8983", x"8982", x"8981", x"8980", x"897f", x"897e", 
    x"897c", x"897b", x"897a", x"8979", x"8978", x"8976", x"8975", x"8974", 
    x"8973", x"8972", x"8971", x"896f", x"896e", x"896d", x"896c", x"896b", 
    x"8969", x"8968", x"8967", x"8966", x"8965", x"8963", x"8962", x"8961", 
    x"8960", x"895f", x"895e", x"895c", x"895b", x"895a", x"8959", x"8958", 
    x"8957", x"8955", x"8954", x"8953", x"8952", x"8951", x"894f", x"894e", 
    x"894d", x"894c", x"894b", x"894a", x"8948", x"8947", x"8946", x"8945", 
    x"8944", x"8943", x"8941", x"8940", x"893f", x"893e", x"893d", x"893c", 
    x"893a", x"8939", x"8938", x"8937", x"8936", x"8934", x"8933", x"8932", 
    x"8931", x"8930", x"892f", x"892d", x"892c", x"892b", x"892a", x"8929", 
    x"8928", x"8926", x"8925", x"8924", x"8923", x"8922", x"8921", x"891f", 
    x"891e", x"891d", x"891c", x"891b", x"891a", x"8919", x"8917", x"8916", 
    x"8915", x"8914", x"8913", x"8912", x"8910", x"890f", x"890e", x"890d", 
    x"890c", x"890b", x"8909", x"8908", x"8907", x"8906", x"8905", x"8904", 
    x"8902", x"8901", x"8900", x"88ff", x"88fe", x"88fd", x"88fc", x"88fa", 
    x"88f9", x"88f8", x"88f7", x"88f6", x"88f5", x"88f3", x"88f2", x"88f1", 
    x"88f0", x"88ef", x"88ee", x"88ed", x"88eb", x"88ea", x"88e9", x"88e8", 
    x"88e7", x"88e6", x"88e4", x"88e3", x"88e2", x"88e1", x"88e0", x"88df", 
    x"88de", x"88dc", x"88db", x"88da", x"88d9", x"88d8", x"88d7", x"88d6", 
    x"88d4", x"88d3", x"88d2", x"88d1", x"88d0", x"88cf", x"88ce", x"88cc", 
    x"88cb", x"88ca", x"88c9", x"88c8", x"88c7", x"88c6", x"88c4", x"88c3", 
    x"88c2", x"88c1", x"88c0", x"88bf", x"88be", x"88bc", x"88bb", x"88ba", 
    x"88b9", x"88b8", x"88b7", x"88b6", x"88b4", x"88b3", x"88b2", x"88b1", 
    x"88b0", x"88af", x"88ae", x"88ac", x"88ab", x"88aa", x"88a9", x"88a8", 
    x"88a7", x"88a6", x"88a4", x"88a3", x"88a2", x"88a1", x"88a0", x"889f", 
    x"889e", x"889d", x"889b", x"889a", x"8899", x"8898", x"8897", x"8896", 
    x"8895", x"8893", x"8892", x"8891", x"8890", x"888f", x"888e", x"888d", 
    x"888c", x"888a", x"8889", x"8888", x"8887", x"8886", x"8885", x"8884", 
    x"8883", x"8881", x"8880", x"887f", x"887e", x"887d", x"887c", x"887b", 
    x"887a", x"8878", x"8877", x"8876", x"8875", x"8874", x"8873", x"8872", 
    x"8871", x"886f", x"886e", x"886d", x"886c", x"886b", x"886a", x"8869", 
    x"8868", x"8867", x"8865", x"8864", x"8863", x"8862", x"8861", x"8860", 
    x"885f", x"885e", x"885c", x"885b", x"885a", x"8859", x"8858", x"8857", 
    x"8856", x"8855", x"8854", x"8852", x"8851", x"8850", x"884f", x"884e", 
    x"884d", x"884c", x"884b", x"884a", x"8848", x"8847", x"8846", x"8845", 
    x"8844", x"8843", x"8842", x"8841", x"8840", x"883e", x"883d", x"883c", 
    x"883b", x"883a", x"8839", x"8838", x"8837", x"8836", x"8834", x"8833", 
    x"8832", x"8831", x"8830", x"882f", x"882e", x"882d", x"882c", x"882a", 
    x"8829", x"8828", x"8827", x"8826", x"8825", x"8824", x"8823", x"8822", 
    x"8821", x"881f", x"881e", x"881d", x"881c", x"881b", x"881a", x"8819", 
    x"8818", x"8817", x"8816", x"8814", x"8813", x"8812", x"8811", x"8810", 
    x"880f", x"880e", x"880d", x"880c", x"880b", x"8809", x"8808", x"8807", 
    x"8806", x"8805", x"8804", x"8803", x"8802", x"8801", x"8800", x"87ff", 
    x"87fd", x"87fc", x"87fb", x"87fa", x"87f9", x"87f8", x"87f7", x"87f6", 
    x"87f5", x"87f4", x"87f3", x"87f1", x"87f0", x"87ef", x"87ee", x"87ed", 
    x"87ec", x"87eb", x"87ea", x"87e9", x"87e8", x"87e7", x"87e6", x"87e4", 
    x"87e3", x"87e2", x"87e1", x"87e0", x"87df", x"87de", x"87dd", x"87dc", 
    x"87db", x"87da", x"87d8", x"87d7", x"87d6", x"87d5", x"87d4", x"87d3", 
    x"87d2", x"87d1", x"87d0", x"87cf", x"87ce", x"87cd", x"87cc", x"87ca", 
    x"87c9", x"87c8", x"87c7", x"87c6", x"87c5", x"87c4", x"87c3", x"87c2", 
    x"87c1", x"87c0", x"87bf", x"87be", x"87bc", x"87bb", x"87ba", x"87b9", 
    x"87b8", x"87b7", x"87b6", x"87b5", x"87b4", x"87b3", x"87b2", x"87b1", 
    x"87b0", x"87ae", x"87ad", x"87ac", x"87ab", x"87aa", x"87a9", x"87a8", 
    x"87a7", x"87a6", x"87a5", x"87a4", x"87a3", x"87a2", x"87a1", x"87a0", 
    x"879e", x"879d", x"879c", x"879b", x"879a", x"8799", x"8798", x"8797", 
    x"8796", x"8795", x"8794", x"8793", x"8792", x"8791", x"8790", x"878e", 
    x"878d", x"878c", x"878b", x"878a", x"8789", x"8788", x"8787", x"8786", 
    x"8785", x"8784", x"8783", x"8782", x"8781", x"8780", x"877f", x"877d", 
    x"877c", x"877b", x"877a", x"8779", x"8778", x"8777", x"8776", x"8775", 
    x"8774", x"8773", x"8772", x"8771", x"8770", x"876f", x"876e", x"876d", 
    x"876c", x"876a", x"8769", x"8768", x"8767", x"8766", x"8765", x"8764", 
    x"8763", x"8762", x"8761", x"8760", x"875f", x"875e", x"875d", x"875c", 
    x"875b", x"875a", x"8759", x"8758", x"8757", x"8755", x"8754", x"8753", 
    x"8752", x"8751", x"8750", x"874f", x"874e", x"874d", x"874c", x"874b", 
    x"874a", x"8749", x"8748", x"8747", x"8746", x"8745", x"8744", x"8743", 
    x"8742", x"8741", x"8740", x"873e", x"873d", x"873c", x"873b", x"873a", 
    x"8739", x"8738", x"8737", x"8736", x"8735", x"8734", x"8733", x"8732", 
    x"8731", x"8730", x"872f", x"872e", x"872d", x"872c", x"872b", x"872a", 
    x"8729", x"8728", x"8727", x"8726", x"8725", x"8723", x"8722", x"8721", 
    x"8720", x"871f", x"871e", x"871d", x"871c", x"871b", x"871a", x"8719", 
    x"8718", x"8717", x"8716", x"8715", x"8714", x"8713", x"8712", x"8711", 
    x"8710", x"870f", x"870e", x"870d", x"870c", x"870b", x"870a", x"8709", 
    x"8708", x"8707", x"8706", x"8705", x"8704", x"8703", x"8702", x"8700", 
    x"86ff", x"86fe", x"86fd", x"86fc", x"86fb", x"86fa", x"86f9", x"86f8", 
    x"86f7", x"86f6", x"86f5", x"86f4", x"86f3", x"86f2", x"86f1", x"86f0", 
    x"86ef", x"86ee", x"86ed", x"86ec", x"86eb", x"86ea", x"86e9", x"86e8", 
    x"86e7", x"86e6", x"86e5", x"86e4", x"86e3", x"86e2", x"86e1", x"86e0", 
    x"86df", x"86de", x"86dd", x"86dc", x"86db", x"86da", x"86d9", x"86d8", 
    x"86d7", x"86d6", x"86d5", x"86d4", x"86d3", x"86d2", x"86d1", x"86d0", 
    x"86cf", x"86ce", x"86cd", x"86cc", x"86cb", x"86ca", x"86c9", x"86c8", 
    x"86c7", x"86c6", x"86c5", x"86c4", x"86c3", x"86c2", x"86c1", x"86c0", 
    x"86bf", x"86bd", x"86bc", x"86bb", x"86ba", x"86b9", x"86b8", x"86b7", 
    x"86b6", x"86b5", x"86b4", x"86b3", x"86b2", x"86b1", x"86b0", x"86af", 
    x"86ae", x"86ad", x"86ac", x"86ab", x"86aa", x"86a9", x"86a8", x"86a7", 
    x"86a6", x"86a5", x"86a4", x"86a3", x"86a2", x"86a1", x"86a0", x"869f", 
    x"869e", x"869d", x"869c", x"869b", x"869a", x"8699", x"8698", x"8697", 
    x"8696", x"8695", x"8695", x"8694", x"8693", x"8692", x"8691", x"8690", 
    x"868f", x"868e", x"868d", x"868c", x"868b", x"868a", x"8689", x"8688", 
    x"8687", x"8686", x"8685", x"8684", x"8683", x"8682", x"8681", x"8680", 
    x"867f", x"867e", x"867d", x"867c", x"867b", x"867a", x"8679", x"8678", 
    x"8677", x"8676", x"8675", x"8674", x"8673", x"8672", x"8671", x"8670", 
    x"866f", x"866e", x"866d", x"866c", x"866b", x"866a", x"8669", x"8668", 
    x"8667", x"8666", x"8665", x"8664", x"8663", x"8662", x"8661", x"8660", 
    x"865f", x"865e", x"865d", x"865c", x"865b", x"865a", x"8659", x"8658", 
    x"8657", x"8656", x"8655", x"8654", x"8654", x"8653", x"8652", x"8651", 
    x"8650", x"864f", x"864e", x"864d", x"864c", x"864b", x"864a", x"8649", 
    x"8648", x"8647", x"8646", x"8645", x"8644", x"8643", x"8642", x"8641", 
    x"8640", x"863f", x"863e", x"863d", x"863c", x"863b", x"863a", x"8639", 
    x"8638", x"8637", x"8636", x"8635", x"8634", x"8633", x"8633", x"8632", 
    x"8631", x"8630", x"862f", x"862e", x"862d", x"862c", x"862b", x"862a", 
    x"8629", x"8628", x"8627", x"8626", x"8625", x"8624", x"8623", x"8622", 
    x"8621", x"8620", x"861f", x"861e", x"861d", x"861c", x"861b", x"861a", 
    x"861a", x"8619", x"8618", x"8617", x"8616", x"8615", x"8614", x"8613", 
    x"8612", x"8611", x"8610", x"860f", x"860e", x"860d", x"860c", x"860b", 
    x"860a", x"8609", x"8608", x"8607", x"8606", x"8605", x"8605", x"8604", 
    x"8603", x"8602", x"8601", x"8600", x"85ff", x"85fe", x"85fd", x"85fc", 
    x"85fb", x"85fa", x"85f9", x"85f8", x"85f7", x"85f6", x"85f5", x"85f4", 
    x"85f3", x"85f2", x"85f2", x"85f1", x"85f0", x"85ef", x"85ee", x"85ed", 
    x"85ec", x"85eb", x"85ea", x"85e9", x"85e8", x"85e7", x"85e6", x"85e5", 
    x"85e4", x"85e3", x"85e2", x"85e2", x"85e1", x"85e0", x"85df", x"85de", 
    x"85dd", x"85dc", x"85db", x"85da", x"85d9", x"85d8", x"85d7", x"85d6", 
    x"85d5", x"85d4", x"85d3", x"85d2", x"85d2", x"85d1", x"85d0", x"85cf", 
    x"85ce", x"85cd", x"85cc", x"85cb", x"85ca", x"85c9", x"85c8", x"85c7", 
    x"85c6", x"85c5", x"85c4", x"85c4", x"85c3", x"85c2", x"85c1", x"85c0", 
    x"85bf", x"85be", x"85bd", x"85bc", x"85bb", x"85ba", x"85b9", x"85b8", 
    x"85b7", x"85b7", x"85b6", x"85b5", x"85b4", x"85b3", x"85b2", x"85b1", 
    x"85b0", x"85af", x"85ae", x"85ad", x"85ac", x"85ab", x"85aa", x"85aa", 
    x"85a9", x"85a8", x"85a7", x"85a6", x"85a5", x"85a4", x"85a3", x"85a2", 
    x"85a1", x"85a0", x"859f", x"859f", x"859e", x"859d", x"859c", x"859b", 
    x"859a", x"8599", x"8598", x"8597", x"8596", x"8595", x"8594", x"8593", 
    x"8593", x"8592", x"8591", x"8590", x"858f", x"858e", x"858d", x"858c", 
    x"858b", x"858a", x"8589", x"8588", x"8588", x"8587", x"8586", x"8585", 
    x"8584", x"8583", x"8582", x"8581", x"8580", x"857f", x"857e", x"857e", 
    x"857d", x"857c", x"857b", x"857a", x"8579", x"8578", x"8577", x"8576", 
    x"8575", x"8574", x"8574", x"8573", x"8572", x"8571", x"8570", x"856f", 
    x"856e", x"856d", x"856c", x"856b", x"856b", x"856a", x"8569", x"8568", 
    x"8567", x"8566", x"8565", x"8564", x"8563", x"8562", x"8561", x"8561", 
    x"8560", x"855f", x"855e", x"855d", x"855c", x"855b", x"855a", x"8559", 
    x"8558", x"8558", x"8557", x"8556", x"8555", x"8554", x"8553", x"8552", 
    x"8551", x"8550", x"8550", x"854f", x"854e", x"854d", x"854c", x"854b", 
    x"854a", x"8549", x"8548", x"8547", x"8547", x"8546", x"8545", x"8544", 
    x"8543", x"8542", x"8541", x"8540", x"853f", x"853f", x"853e", x"853d", 
    x"853c", x"853b", x"853a", x"8539", x"8538", x"8537", x"8537", x"8536", 
    x"8535", x"8534", x"8533", x"8532", x"8531", x"8530", x"852f", x"852f", 
    x"852e", x"852d", x"852c", x"852b", x"852a", x"8529", x"8528", x"8528", 
    x"8527", x"8526", x"8525", x"8524", x"8523", x"8522", x"8521", x"8520", 
    x"8520", x"851f", x"851e", x"851d", x"851c", x"851b", x"851a", x"8519", 
    x"8519", x"8518", x"8517", x"8516", x"8515", x"8514", x"8513", x"8512", 
    x"8512", x"8511", x"8510", x"850f", x"850e", x"850d", x"850c", x"850b", 
    x"850b", x"850a", x"8509", x"8508", x"8507", x"8506", x"8505", x"8504", 
    x"8504", x"8503", x"8502", x"8501", x"8500", x"84ff", x"84fe", x"84fe", 
    x"84fd", x"84fc", x"84fb", x"84fa", x"84f9", x"84f8", x"84f7", x"84f7", 
    x"84f6", x"84f5", x"84f4", x"84f3", x"84f2", x"84f1", x"84f1", x"84f0", 
    x"84ef", x"84ee", x"84ed", x"84ec", x"84eb", x"84ea", x"84ea", x"84e9", 
    x"84e8", x"84e7", x"84e6", x"84e5", x"84e4", x"84e4", x"84e3", x"84e2", 
    x"84e1", x"84e0", x"84df", x"84de", x"84de", x"84dd", x"84dc", x"84db", 
    x"84da", x"84d9", x"84d8", x"84d8", x"84d7", x"84d6", x"84d5", x"84d4", 
    x"84d3", x"84d2", x"84d2", x"84d1", x"84d0", x"84cf", x"84ce", x"84cd", 
    x"84cd", x"84cc", x"84cb", x"84ca", x"84c9", x"84c8", x"84c7", x"84c7", 
    x"84c6", x"84c5", x"84c4", x"84c3", x"84c2", x"84c1", x"84c1", x"84c0", 
    x"84bf", x"84be", x"84bd", x"84bc", x"84bc", x"84bb", x"84ba", x"84b9", 
    x"84b8", x"84b7", x"84b6", x"84b6", x"84b5", x"84b4", x"84b3", x"84b2", 
    x"84b1", x"84b1", x"84b0", x"84af", x"84ae", x"84ad", x"84ac", x"84ac", 
    x"84ab", x"84aa", x"84a9", x"84a8", x"84a7", x"84a6", x"84a6", x"84a5", 
    x"84a4", x"84a3", x"84a2", x"84a1", x"84a1", x"84a0", x"849f", x"849e", 
    x"849d", x"849c", x"849c", x"849b", x"849a", x"8499", x"8498", x"8497", 
    x"8497", x"8496", x"8495", x"8494", x"8493", x"8492", x"8492", x"8491", 
    x"8490", x"848f", x"848e", x"848d", x"848d", x"848c", x"848b", x"848a", 
    x"8489", x"8488", x"8488", x"8487", x"8486", x"8485", x"8484", x"8483", 
    x"8483", x"8482", x"8481", x"8480", x"847f", x"847f", x"847e", x"847d", 
    x"847c", x"847b", x"847a", x"847a", x"8479", x"8478", x"8477", x"8476", 
    x"8475", x"8475", x"8474", x"8473", x"8472", x"8471", x"8471", x"8470", 
    x"846f", x"846e", x"846d", x"846c", x"846c", x"846b", x"846a", x"8469", 
    x"8468", x"8468", x"8467", x"8466", x"8465", x"8464", x"8463", x"8463", 
    x"8462", x"8461", x"8460", x"845f", x"845f", x"845e", x"845d", x"845c", 
    x"845b", x"845b", x"845a", x"8459", x"8458", x"8457", x"8456", x"8456", 
    x"8455", x"8454", x"8453", x"8452", x"8452", x"8451", x"8450", x"844f", 
    x"844e", x"844e", x"844d", x"844c", x"844b", x"844a", x"844a", x"8449", 
    x"8448", x"8447", x"8446", x"8446", x"8445", x"8444", x"8443", x"8442", 
    x"8441", x"8441", x"8440", x"843f", x"843e", x"843d", x"843d", x"843c", 
    x"843b", x"843a", x"8439", x"8439", x"8438", x"8437", x"8436", x"8435", 
    x"8435", x"8434", x"8433", x"8432", x"8431", x"8431", x"8430", x"842f", 
    x"842e", x"842e", x"842d", x"842c", x"842b", x"842a", x"842a", x"8429", 
    x"8428", x"8427", x"8426", x"8426", x"8425", x"8424", x"8423", x"8422", 
    x"8422", x"8421", x"8420", x"841f", x"841e", x"841e", x"841d", x"841c", 
    x"841b", x"841a", x"841a", x"8419", x"8418", x"8417", x"8417", x"8416", 
    x"8415", x"8414", x"8413", x"8413", x"8412", x"8411", x"8410", x"840f", 
    x"840f", x"840e", x"840d", x"840c", x"840c", x"840b", x"840a", x"8409", 
    x"8408", x"8408", x"8407", x"8406", x"8405", x"8405", x"8404", x"8403", 
    x"8402", x"8401", x"8401", x"8400", x"83ff", x"83fe", x"83fe", x"83fd", 
    x"83fc", x"83fb", x"83fa", x"83fa", x"83f9", x"83f8", x"83f7", x"83f7", 
    x"83f6", x"83f5", x"83f4", x"83f3", x"83f3", x"83f2", x"83f1", x"83f0", 
    x"83f0", x"83ef", x"83ee", x"83ed", x"83ec", x"83ec", x"83eb", x"83ea", 
    x"83e9", x"83e9", x"83e8", x"83e7", x"83e6", x"83e6", x"83e5", x"83e4", 
    x"83e3", x"83e2", x"83e2", x"83e1", x"83e0", x"83df", x"83df", x"83de", 
    x"83dd", x"83dc", x"83dc", x"83db", x"83da", x"83d9", x"83d9", x"83d8", 
    x"83d7", x"83d6", x"83d5", x"83d5", x"83d4", x"83d3", x"83d2", x"83d2", 
    x"83d1", x"83d0", x"83cf", x"83cf", x"83ce", x"83cd", x"83cc", x"83cc", 
    x"83cb", x"83ca", x"83c9", x"83c9", x"83c8", x"83c7", x"83c6", x"83c6", 
    x"83c5", x"83c4", x"83c3", x"83c2", x"83c2", x"83c1", x"83c0", x"83bf", 
    x"83bf", x"83be", x"83bd", x"83bc", x"83bc", x"83bb", x"83ba", x"83b9", 
    x"83b9", x"83b8", x"83b7", x"83b6", x"83b6", x"83b5", x"83b4", x"83b3", 
    x"83b3", x"83b2", x"83b1", x"83b0", x"83b0", x"83af", x"83ae", x"83ad", 
    x"83ad", x"83ac", x"83ab", x"83aa", x"83aa", x"83a9", x"83a8", x"83a7", 
    x"83a7", x"83a6", x"83a5", x"83a4", x"83a4", x"83a3", x"83a2", x"83a2", 
    x"83a1", x"83a0", x"839f", x"839f", x"839e", x"839d", x"839c", x"839c", 
    x"839b", x"839a", x"8399", x"8399", x"8398", x"8397", x"8396", x"8396", 
    x"8395", x"8394", x"8393", x"8393", x"8392", x"8391", x"8391", x"8390", 
    x"838f", x"838e", x"838e", x"838d", x"838c", x"838b", x"838b", x"838a", 
    x"8389", x"8388", x"8388", x"8387", x"8386", x"8386", x"8385", x"8384", 
    x"8383", x"8383", x"8382", x"8381", x"8380", x"8380", x"837f", x"837e", 
    x"837d", x"837d", x"837c", x"837b", x"837b", x"837a", x"8379", x"8378", 
    x"8378", x"8377", x"8376", x"8376", x"8375", x"8374", x"8373", x"8373", 
    x"8372", x"8371", x"8370", x"8370", x"836f", x"836e", x"836e", x"836d", 
    x"836c", x"836b", x"836b", x"836a", x"8369", x"8368", x"8368", x"8367", 
    x"8366", x"8366", x"8365", x"8364", x"8363", x"8363", x"8362", x"8361", 
    x"8361", x"8360", x"835f", x"835e", x"835e", x"835d", x"835c", x"835c", 
    x"835b", x"835a", x"8359", x"8359", x"8358", x"8357", x"8357", x"8356", 
    x"8355", x"8354", x"8354", x"8353", x"8352", x"8352", x"8351", x"8350", 
    x"834f", x"834f", x"834e", x"834d", x"834d", x"834c", x"834b", x"834b", 
    x"834a", x"8349", x"8348", x"8348", x"8347", x"8346", x"8346", x"8345", 
    x"8344", x"8343", x"8343", x"8342", x"8341", x"8341", x"8340", x"833f", 
    x"833f", x"833e", x"833d", x"833c", x"833c", x"833b", x"833a", x"833a", 
    x"8339", x"8338", x"8338", x"8337", x"8336", x"8335", x"8335", x"8334", 
    x"8333", x"8333", x"8332", x"8331", x"8331", x"8330", x"832f", x"832e", 
    x"832e", x"832d", x"832c", x"832c", x"832b", x"832a", x"832a", x"8329", 
    x"8328", x"8328", x"8327", x"8326", x"8325", x"8325", x"8324", x"8323", 
    x"8323", x"8322", x"8321", x"8321", x"8320", x"831f", x"831f", x"831e", 
    x"831d", x"831c", x"831c", x"831b", x"831a", x"831a", x"8319", x"8318", 
    x"8318", x"8317", x"8316", x"8316", x"8315", x"8314", x"8314", x"8313", 
    x"8312", x"8312", x"8311", x"8310", x"830f", x"830f", x"830e", x"830d", 
    x"830d", x"830c", x"830b", x"830b", x"830a", x"8309", x"8309", x"8308", 
    x"8307", x"8307", x"8306", x"8305", x"8305", x"8304", x"8303", x"8303", 
    x"8302", x"8301", x"8301", x"8300", x"82ff", x"82fe", x"82fe", x"82fd", 
    x"82fc", x"82fc", x"82fb", x"82fa", x"82fa", x"82f9", x"82f8", x"82f8", 
    x"82f7", x"82f6", x"82f6", x"82f5", x"82f4", x"82f4", x"82f3", x"82f2", 
    x"82f2", x"82f1", x"82f0", x"82f0", x"82ef", x"82ee", x"82ee", x"82ed", 
    x"82ec", x"82ec", x"82eb", x"82ea", x"82ea", x"82e9", x"82e8", x"82e8", 
    x"82e7", x"82e6", x"82e6", x"82e5", x"82e4", x"82e4", x"82e3", x"82e2", 
    x"82e2", x"82e1", x"82e0", x"82e0", x"82df", x"82de", x"82de", x"82dd", 
    x"82dc", x"82dc", x"82db", x"82da", x"82da", x"82d9", x"82d8", x"82d8", 
    x"82d7", x"82d7", x"82d6", x"82d5", x"82d5", x"82d4", x"82d3", x"82d3", 
    x"82d2", x"82d1", x"82d1", x"82d0", x"82cf", x"82cf", x"82ce", x"82cd", 
    x"82cd", x"82cc", x"82cb", x"82cb", x"82ca", x"82c9", x"82c9", x"82c8", 
    x"82c7", x"82c7", x"82c6", x"82c6", x"82c5", x"82c4", x"82c4", x"82c3", 
    x"82c2", x"82c2", x"82c1", x"82c0", x"82c0", x"82bf", x"82be", x"82be", 
    x"82bd", x"82bc", x"82bc", x"82bb", x"82bb", x"82ba", x"82b9", x"82b9", 
    x"82b8", x"82b7", x"82b7", x"82b6", x"82b5", x"82b5", x"82b4", x"82b3", 
    x"82b3", x"82b2", x"82b2", x"82b1", x"82b0", x"82b0", x"82af", x"82ae", 
    x"82ae", x"82ad", x"82ac", x"82ac", x"82ab", x"82aa", x"82aa", x"82a9", 
    x"82a9", x"82a8", x"82a7", x"82a7", x"82a6", x"82a5", x"82a5", x"82a4", 
    x"82a4", x"82a3", x"82a2", x"82a2", x"82a1", x"82a0", x"82a0", x"829f", 
    x"829e", x"829e", x"829d", x"829d", x"829c", x"829b", x"829b", x"829a", 
    x"8299", x"8299", x"8298", x"8298", x"8297", x"8296", x"8296", x"8295", 
    x"8294", x"8294", x"8293", x"8292", x"8292", x"8291", x"8291", x"8290", 
    x"828f", x"828f", x"828e", x"828d", x"828d", x"828c", x"828c", x"828b", 
    x"828a", x"828a", x"8289", x"8289", x"8288", x"8287", x"8287", x"8286", 
    x"8285", x"8285", x"8284", x"8284", x"8283", x"8282", x"8282", x"8281", 
    x"8280", x"8280", x"827f", x"827f", x"827e", x"827d", x"827d", x"827c", 
    x"827c", x"827b", x"827a", x"827a", x"8279", x"8278", x"8278", x"8277", 
    x"8277", x"8276", x"8275", x"8275", x"8274", x"8274", x"8273", x"8272", 
    x"8272", x"8271", x"8270", x"8270", x"826f", x"826f", x"826e", x"826d", 
    x"826d", x"826c", x"826c", x"826b", x"826a", x"826a", x"8269", x"8269", 
    x"8268", x"8267", x"8267", x"8266", x"8266", x"8265", x"8264", x"8264", 
    x"8263", x"8263", x"8262", x"8261", x"8261", x"8260", x"8260", x"825f", 
    x"825e", x"825e", x"825d", x"825d", x"825c", x"825b", x"825b", x"825a", 
    x"825a", x"8259", x"8258", x"8258", x"8257", x"8257", x"8256", x"8255", 
    x"8255", x"8254", x"8254", x"8253", x"8252", x"8252", x"8251", x"8251", 
    x"8250", x"824f", x"824f", x"824e", x"824e", x"824d", x"824c", x"824c", 
    x"824b", x"824b", x"824a", x"8249", x"8249", x"8248", x"8248", x"8247", 
    x"8247", x"8246", x"8245", x"8245", x"8244", x"8244", x"8243", x"8242", 
    x"8242", x"8241", x"8241", x"8240", x"823f", x"823f", x"823e", x"823e", 
    x"823d", x"823d", x"823c", x"823b", x"823b", x"823a", x"823a", x"8239", 
    x"8238", x"8238", x"8237", x"8237", x"8236", x"8236", x"8235", x"8234", 
    x"8234", x"8233", x"8233", x"8232", x"8232", x"8231", x"8230", x"8230", 
    x"822f", x"822f", x"822e", x"822d", x"822d", x"822c", x"822c", x"822b", 
    x"822b", x"822a", x"8229", x"8229", x"8228", x"8228", x"8227", x"8227", 
    x"8226", x"8225", x"8225", x"8224", x"8224", x"8223", x"8223", x"8222", 
    x"8221", x"8221", x"8220", x"8220", x"821f", x"821f", x"821e", x"821d", 
    x"821d", x"821c", x"821c", x"821b", x"821b", x"821a", x"8219", x"8219", 
    x"8218", x"8218", x"8217", x"8217", x"8216", x"8216", x"8215", x"8214", 
    x"8214", x"8213", x"8213", x"8212", x"8212", x"8211", x"8210", x"8210", 
    x"820f", x"820f", x"820e", x"820e", x"820d", x"820d", x"820c", x"820b", 
    x"820b", x"820a", x"820a", x"8209", x"8209", x"8208", x"8208", x"8207", 
    x"8206", x"8206", x"8205", x"8205", x"8204", x"8204", x"8203", x"8203", 
    x"8202", x"8201", x"8201", x"8200", x"8200", x"81ff", x"81ff", x"81fe", 
    x"81fe", x"81fd", x"81fc", x"81fc", x"81fb", x"81fb", x"81fa", x"81fa", 
    x"81f9", x"81f9", x"81f8", x"81f7", x"81f7", x"81f6", x"81f6", x"81f5", 
    x"81f5", x"81f4", x"81f4", x"81f3", x"81f3", x"81f2", x"81f1", x"81f1", 
    x"81f0", x"81f0", x"81ef", x"81ef", x"81ee", x"81ee", x"81ed", x"81ed", 
    x"81ec", x"81eb", x"81eb", x"81ea", x"81ea", x"81e9", x"81e9", x"81e8", 
    x"81e8", x"81e7", x"81e7", x"81e6", x"81e6", x"81e5", x"81e4", x"81e4", 
    x"81e3", x"81e3", x"81e2", x"81e2", x"81e1", x"81e1", x"81e0", x"81e0", 
    x"81df", x"81df", x"81de", x"81de", x"81dd", x"81dc", x"81dc", x"81db", 
    x"81db", x"81da", x"81da", x"81d9", x"81d9", x"81d8", x"81d8", x"81d7", 
    x"81d7", x"81d6", x"81d6", x"81d5", x"81d4", x"81d4", x"81d3", x"81d3", 
    x"81d2", x"81d2", x"81d1", x"81d1", x"81d0", x"81d0", x"81cf", x"81cf", 
    x"81ce", x"81ce", x"81cd", x"81cd", x"81cc", x"81cc", x"81cb", x"81ca", 
    x"81ca", x"81c9", x"81c9", x"81c8", x"81c8", x"81c7", x"81c7", x"81c6", 
    x"81c6", x"81c5", x"81c5", x"81c4", x"81c4", x"81c3", x"81c3", x"81c2", 
    x"81c2", x"81c1", x"81c1", x"81c0", x"81c0", x"81bf", x"81bf", x"81be", 
    x"81be", x"81bd", x"81bc", x"81bc", x"81bb", x"81bb", x"81ba", x"81ba", 
    x"81b9", x"81b9", x"81b8", x"81b8", x"81b7", x"81b7", x"81b6", x"81b6", 
    x"81b5", x"81b5", x"81b4", x"81b4", x"81b3", x"81b3", x"81b2", x"81b2", 
    x"81b1", x"81b1", x"81b0", x"81b0", x"81af", x"81af", x"81ae", x"81ae", 
    x"81ad", x"81ad", x"81ac", x"81ac", x"81ab", x"81ab", x"81aa", x"81aa", 
    x"81a9", x"81a9", x"81a8", x"81a8", x"81a7", x"81a7", x"81a6", x"81a6", 
    x"81a5", x"81a5", x"81a4", x"81a4", x"81a3", x"81a3", x"81a2", x"81a2", 
    x"81a1", x"81a1", x"81a0", x"81a0", x"819f", x"819f", x"819e", x"819e", 
    x"819d", x"819d", x"819c", x"819c", x"819b", x"819b", x"819a", x"819a", 
    x"8199", x"8199", x"8198", x"8198", x"8197", x"8197", x"8196", x"8196", 
    x"8195", x"8195", x"8194", x"8194", x"8193", x"8193", x"8192", x"8192", 
    x"8191", x"8191", x"8190", x"8190", x"818f", x"818f", x"818e", x"818e", 
    x"818d", x"818d", x"818c", x"818c", x"818b", x"818b", x"818a", x"818a", 
    x"8189", x"8189", x"8189", x"8188", x"8188", x"8187", x"8187", x"8186", 
    x"8186", x"8185", x"8185", x"8184", x"8184", x"8183", x"8183", x"8182", 
    x"8182", x"8181", x"8181", x"8180", x"8180", x"817f", x"817f", x"817e", 
    x"817e", x"817d", x"817d", x"817d", x"817c", x"817c", x"817b", x"817b", 
    x"817a", x"817a", x"8179", x"8179", x"8178", x"8178", x"8177", x"8177", 
    x"8176", x"8176", x"8175", x"8175", x"8174", x"8174", x"8173", x"8173", 
    x"8173", x"8172", x"8172", x"8171", x"8171", x"8170", x"8170", x"816f", 
    x"816f", x"816e", x"816e", x"816d", x"816d", x"816c", x"816c", x"816c", 
    x"816b", x"816b", x"816a", x"816a", x"8169", x"8169", x"8168", x"8168", 
    x"8167", x"8167", x"8166", x"8166", x"8165", x"8165", x"8165", x"8164", 
    x"8164", x"8163", x"8163", x"8162", x"8162", x"8161", x"8161", x"8160", 
    x"8160", x"8160", x"815f", x"815f", x"815e", x"815e", x"815d", x"815d", 
    x"815c", x"815c", x"815b", x"815b", x"815a", x"815a", x"815a", x"8159", 
    x"8159", x"8158", x"8158", x"8157", x"8157", x"8156", x"8156", x"8156", 
    x"8155", x"8155", x"8154", x"8154", x"8153", x"8153", x"8152", x"8152", 
    x"8151", x"8151", x"8151", x"8150", x"8150", x"814f", x"814f", x"814e", 
    x"814e", x"814d", x"814d", x"814d", x"814c", x"814c", x"814b", x"814b", 
    x"814a", x"814a", x"8149", x"8149", x"8149", x"8148", x"8148", x"8147", 
    x"8147", x"8146", x"8146", x"8145", x"8145", x"8145", x"8144", x"8144", 
    x"8143", x"8143", x"8142", x"8142", x"8141", x"8141", x"8141", x"8140", 
    x"8140", x"813f", x"813f", x"813e", x"813e", x"813e", x"813d", x"813d", 
    x"813c", x"813c", x"813b", x"813b", x"813b", x"813a", x"813a", x"8139", 
    x"8139", x"8138", x"8138", x"8137", x"8137", x"8137", x"8136", x"8136", 
    x"8135", x"8135", x"8134", x"8134", x"8134", x"8133", x"8133", x"8132", 
    x"8132", x"8131", x"8131", x"8131", x"8130", x"8130", x"812f", x"812f", 
    x"812e", x"812e", x"812e", x"812d", x"812d", x"812c", x"812c", x"812c", 
    x"812b", x"812b", x"812a", x"812a", x"8129", x"8129", x"8129", x"8128", 
    x"8128", x"8127", x"8127", x"8126", x"8126", x"8126", x"8125", x"8125", 
    x"8124", x"8124", x"8124", x"8123", x"8123", x"8122", x"8122", x"8121", 
    x"8121", x"8121", x"8120", x"8120", x"811f", x"811f", x"811f", x"811e", 
    x"811e", x"811d", x"811d", x"811c", x"811c", x"811c", x"811b", x"811b", 
    x"811a", x"811a", x"811a", x"8119", x"8119", x"8118", x"8118", x"8118", 
    x"8117", x"8117", x"8116", x"8116", x"8116", x"8115", x"8115", x"8114", 
    x"8114", x"8113", x"8113", x"8113", x"8112", x"8112", x"8111", x"8111", 
    x"8111", x"8110", x"8110", x"810f", x"810f", x"810f", x"810e", x"810e", 
    x"810d", x"810d", x"810d", x"810c", x"810c", x"810b", x"810b", x"810b", 
    x"810a", x"810a", x"8109", x"8109", x"8109", x"8108", x"8108", x"8107", 
    x"8107", x"8107", x"8106", x"8106", x"8105", x"8105", x"8105", x"8104", 
    x"8104", x"8103", x"8103", x"8103", x"8102", x"8102", x"8102", x"8101", 
    x"8101", x"8100", x"8100", x"8100", x"80ff", x"80ff", x"80fe", x"80fe", 
    x"80fe", x"80fd", x"80fd", x"80fc", x"80fc", x"80fc", x"80fb", x"80fb", 
    x"80fb", x"80fa", x"80fa", x"80f9", x"80f9", x"80f9", x"80f8", x"80f8", 
    x"80f7", x"80f7", x"80f7", x"80f6", x"80f6", x"80f6", x"80f5", x"80f5", 
    x"80f4", x"80f4", x"80f4", x"80f3", x"80f3", x"80f2", x"80f2", x"80f2", 
    x"80f1", x"80f1", x"80f1", x"80f0", x"80f0", x"80ef", x"80ef", x"80ef", 
    x"80ee", x"80ee", x"80ee", x"80ed", x"80ed", x"80ec", x"80ec", x"80ec", 
    x"80eb", x"80eb", x"80eb", x"80ea", x"80ea", x"80e9", x"80e9", x"80e9", 
    x"80e8", x"80e8", x"80e8", x"80e7", x"80e7", x"80e6", x"80e6", x"80e6", 
    x"80e5", x"80e5", x"80e5", x"80e4", x"80e4", x"80e3", x"80e3", x"80e3", 
    x"80e2", x"80e2", x"80e2", x"80e1", x"80e1", x"80e1", x"80e0", x"80e0", 
    x"80df", x"80df", x"80df", x"80de", x"80de", x"80de", x"80dd", x"80dd", 
    x"80dd", x"80dc", x"80dc", x"80db", x"80db", x"80db", x"80da", x"80da", 
    x"80da", x"80d9", x"80d9", x"80d9", x"80d8", x"80d8", x"80d7", x"80d7", 
    x"80d7", x"80d6", x"80d6", x"80d6", x"80d5", x"80d5", x"80d5", x"80d4", 
    x"80d4", x"80d4", x"80d3", x"80d3", x"80d2", x"80d2", x"80d2", x"80d1", 
    x"80d1", x"80d1", x"80d0", x"80d0", x"80d0", x"80cf", x"80cf", x"80cf", 
    x"80ce", x"80ce", x"80ce", x"80cd", x"80cd", x"80cc", x"80cc", x"80cc", 
    x"80cb", x"80cb", x"80cb", x"80ca", x"80ca", x"80ca", x"80c9", x"80c9", 
    x"80c9", x"80c8", x"80c8", x"80c8", x"80c7", x"80c7", x"80c7", x"80c6", 
    x"80c6", x"80c6", x"80c5", x"80c5", x"80c5", x"80c4", x"80c4", x"80c3", 
    x"80c3", x"80c3", x"80c2", x"80c2", x"80c2", x"80c1", x"80c1", x"80c1", 
    x"80c0", x"80c0", x"80c0", x"80bf", x"80bf", x"80bf", x"80be", x"80be", 
    x"80be", x"80bd", x"80bd", x"80bd", x"80bc", x"80bc", x"80bc", x"80bb", 
    x"80bb", x"80bb", x"80ba", x"80ba", x"80ba", x"80b9", x"80b9", x"80b9", 
    x"80b8", x"80b8", x"80b8", x"80b7", x"80b7", x"80b7", x"80b6", x"80b6", 
    x"80b6", x"80b5", x"80b5", x"80b5", x"80b4", x"80b4", x"80b4", x"80b3", 
    x"80b3", x"80b3", x"80b2", x"80b2", x"80b2", x"80b1", x"80b1", x"80b1", 
    x"80b0", x"80b0", x"80b0", x"80b0", x"80af", x"80af", x"80af", x"80ae", 
    x"80ae", x"80ae", x"80ad", x"80ad", x"80ad", x"80ac", x"80ac", x"80ac", 
    x"80ab", x"80ab", x"80ab", x"80aa", x"80aa", x"80aa", x"80a9", x"80a9", 
    x"80a9", x"80a8", x"80a8", x"80a8", x"80a8", x"80a7", x"80a7", x"80a7", 
    x"80a6", x"80a6", x"80a6", x"80a5", x"80a5", x"80a5", x"80a4", x"80a4", 
    x"80a4", x"80a3", x"80a3", x"80a3", x"80a2", x"80a2", x"80a2", x"80a2", 
    x"80a1", x"80a1", x"80a1", x"80a0", x"80a0", x"80a0", x"809f", x"809f", 
    x"809f", x"809e", x"809e", x"809e", x"809e", x"809d", x"809d", x"809d", 
    x"809c", x"809c", x"809c", x"809b", x"809b", x"809b", x"809b", x"809a", 
    x"809a", x"809a", x"8099", x"8099", x"8099", x"8098", x"8098", x"8098", 
    x"8097", x"8097", x"8097", x"8097", x"8096", x"8096", x"8096", x"8095", 
    x"8095", x"8095", x"8094", x"8094", x"8094", x"8094", x"8093", x"8093", 
    x"8093", x"8092", x"8092", x"8092", x"8092", x"8091", x"8091", x"8091", 
    x"8090", x"8090", x"8090", x"808f", x"808f", x"808f", x"808f", x"808e", 
    x"808e", x"808e", x"808d", x"808d", x"808d", x"808d", x"808c", x"808c", 
    x"808c", x"808b", x"808b", x"808b", x"808b", x"808a", x"808a", x"808a", 
    x"8089", x"8089", x"8089", x"8089", x"8088", x"8088", x"8088", x"8087", 
    x"8087", x"8087", x"8087", x"8086", x"8086", x"8086", x"8085", x"8085", 
    x"8085", x"8085", x"8084", x"8084", x"8084", x"8083", x"8083", x"8083", 
    x"8083", x"8082", x"8082", x"8082", x"8081", x"8081", x"8081", x"8081", 
    x"8080", x"8080", x"8080", x"8080", x"807f", x"807f", x"807f", x"807e", 
    x"807e", x"807e", x"807e", x"807d", x"807d", x"807d", x"807d", x"807c", 
    x"807c", x"807c", x"807b", x"807b", x"807b", x"807b", x"807a", x"807a", 
    x"807a", x"807a", x"8079", x"8079", x"8079", x"8078", x"8078", x"8078", 
    x"8078", x"8077", x"8077", x"8077", x"8077", x"8076", x"8076", x"8076", 
    x"8076", x"8075", x"8075", x"8075", x"8074", x"8074", x"8074", x"8074", 
    x"8073", x"8073", x"8073", x"8073", x"8072", x"8072", x"8072", x"8072", 
    x"8071", x"8071", x"8071", x"8071", x"8070", x"8070", x"8070", x"8070", 
    x"806f", x"806f", x"806f", x"806f", x"806e", x"806e", x"806e", x"806d", 
    x"806d", x"806d", x"806d", x"806c", x"806c", x"806c", x"806c", x"806b", 
    x"806b", x"806b", x"806b", x"806a", x"806a", x"806a", x"806a", x"8069", 
    x"8069", x"8069", x"8069", x"8068", x"8068", x"8068", x"8068", x"8067", 
    x"8067", x"8067", x"8067", x"8066", x"8066", x"8066", x"8066", x"8065", 
    x"8065", x"8065", x"8065", x"8064", x"8064", x"8064", x"8064", x"8064", 
    x"8063", x"8063", x"8063", x"8063", x"8062", x"8062", x"8062", x"8062", 
    x"8061", x"8061", x"8061", x"8061", x"8060", x"8060", x"8060", x"8060", 
    x"805f", x"805f", x"805f", x"805f", x"805e", x"805e", x"805e", x"805e", 
    x"805e", x"805d", x"805d", x"805d", x"805d", x"805c", x"805c", x"805c", 
    x"805c", x"805b", x"805b", x"805b", x"805b", x"805a", x"805a", x"805a", 
    x"805a", x"805a", x"8059", x"8059", x"8059", x"8059", x"8058", x"8058", 
    x"8058", x"8058", x"8057", x"8057", x"8057", x"8057", x"8057", x"8056", 
    x"8056", x"8056", x"8056", x"8055", x"8055", x"8055", x"8055", x"8055", 
    x"8054", x"8054", x"8054", x"8054", x"8053", x"8053", x"8053", x"8053", 
    x"8053", x"8052", x"8052", x"8052", x"8052", x"8051", x"8051", x"8051", 
    x"8051", x"8051", x"8050", x"8050", x"8050", x"8050", x"804f", x"804f", 
    x"804f", x"804f", x"804f", x"804e", x"804e", x"804e", x"804e", x"804e", 
    x"804d", x"804d", x"804d", x"804d", x"804c", x"804c", x"804c", x"804c", 
    x"804c", x"804b", x"804b", x"804b", x"804b", x"804b", x"804a", x"804a", 
    x"804a", x"804a", x"804a", x"8049", x"8049", x"8049", x"8049", x"8048", 
    x"8048", x"8048", x"8048", x"8048", x"8047", x"8047", x"8047", x"8047", 
    x"8047", x"8046", x"8046", x"8046", x"8046", x"8046", x"8045", x"8045", 
    x"8045", x"8045", x"8045", x"8044", x"8044", x"8044", x"8044", x"8044", 
    x"8043", x"8043", x"8043", x"8043", x"8043", x"8042", x"8042", x"8042", 
    x"8042", x"8042", x"8041", x"8041", x"8041", x"8041", x"8041", x"8040", 
    x"8040", x"8040", x"8040", x"8040", x"803f", x"803f", x"803f", x"803f", 
    x"803f", x"803e", x"803e", x"803e", x"803e", x"803e", x"803e", x"803d", 
    x"803d", x"803d", x"803d", x"803d", x"803c", x"803c", x"803c", x"803c", 
    x"803c", x"803b", x"803b", x"803b", x"803b", x"803b", x"803a", x"803a", 
    x"803a", x"803a", x"803a", x"803a", x"8039", x"8039", x"8039", x"8039", 
    x"8039", x"8038", x"8038", x"8038", x"8038", x"8038", x"8038", x"8037", 
    x"8037", x"8037", x"8037", x"8037", x"8036", x"8036", x"8036", x"8036", 
    x"8036", x"8036", x"8035", x"8035", x"8035", x"8035", x"8035", x"8035", 
    x"8034", x"8034", x"8034", x"8034", x"8034", x"8033", x"8033", x"8033", 
    x"8033", x"8033", x"8033", x"8032", x"8032", x"8032", x"8032", x"8032", 
    x"8032", x"8031", x"8031", x"8031", x"8031", x"8031", x"8031", x"8030", 
    x"8030", x"8030", x"8030", x"8030", x"8030", x"802f", x"802f", x"802f", 
    x"802f", x"802f", x"802f", x"802e", x"802e", x"802e", x"802e", x"802e", 
    x"802e", x"802d", x"802d", x"802d", x"802d", x"802d", x"802d", x"802c", 
    x"802c", x"802c", x"802c", x"802c", x"802c", x"802b", x"802b", x"802b", 
    x"802b", x"802b", x"802b", x"802a", x"802a", x"802a", x"802a", x"802a", 
    x"802a", x"802a", x"8029", x"8029", x"8029", x"8029", x"8029", x"8029", 
    x"8028", x"8028", x"8028", x"8028", x"8028", x"8028", x"8028", x"8027", 
    x"8027", x"8027", x"8027", x"8027", x"8027", x"8026", x"8026", x"8026", 
    x"8026", x"8026", x"8026", x"8026", x"8025", x"8025", x"8025", x"8025", 
    x"8025", x"8025", x"8025", x"8024", x"8024", x"8024", x"8024", x"8024", 
    x"8024", x"8024", x"8023", x"8023", x"8023", x"8023", x"8023", x"8023", 
    x"8023", x"8022", x"8022", x"8022", x"8022", x"8022", x"8022", x"8022", 
    x"8021", x"8021", x"8021", x"8021", x"8021", x"8021", x"8021", x"8020", 
    x"8020", x"8020", x"8020", x"8020", x"8020", x"8020", x"801f", x"801f", 
    x"801f", x"801f", x"801f", x"801f", x"801f", x"801f", x"801e", x"801e", 
    x"801e", x"801e", x"801e", x"801e", x"801e", x"801d", x"801d", x"801d", 
    x"801d", x"801d", x"801d", x"801d", x"801d", x"801c", x"801c", x"801c", 
    x"801c", x"801c", x"801c", x"801c", x"801c", x"801b", x"801b", x"801b", 
    x"801b", x"801b", x"801b", x"801b", x"801b", x"801a", x"801a", x"801a", 
    x"801a", x"801a", x"801a", x"801a", x"801a", x"8019", x"8019", x"8019", 
    x"8019", x"8019", x"8019", x"8019", x"8019", x"8018", x"8018", x"8018", 
    x"8018", x"8018", x"8018", x"8018", x"8018", x"8018", x"8017", x"8017", 
    x"8017", x"8017", x"8017", x"8017", x"8017", x"8017", x"8017", x"8016", 
    x"8016", x"8016", x"8016", x"8016", x"8016", x"8016", x"8016", x"8016", 
    x"8015", x"8015", x"8015", x"8015", x"8015", x"8015", x"8015", x"8015", 
    x"8015", x"8014", x"8014", x"8014", x"8014", x"8014", x"8014", x"8014", 
    x"8014", x"8014", x"8013", x"8013", x"8013", x"8013", x"8013", x"8013", 
    x"8013", x"8013", x"8013", x"8013", x"8012", x"8012", x"8012", x"8012", 
    x"8012", x"8012", x"8012", x"8012", x"8012", x"8011", x"8011", x"8011", 
    x"8011", x"8011", x"8011", x"8011", x"8011", x"8011", x"8011", x"8011", 
    x"8010", x"8010", x"8010", x"8010", x"8010", x"8010", x"8010", x"8010", 
    x"8010", x"8010", x"800f", x"800f", x"800f", x"800f", x"800f", x"800f", 
    x"800f", x"800f", x"800f", x"800f", x"800f", x"800e", x"800e", x"800e", 
    x"800e", x"800e", x"800e", x"800e", x"800e", x"800e", x"800e", x"800e", 
    x"800d", x"800d", x"800d", x"800d", x"800d", x"800d", x"800d", x"800d", 
    x"800d", x"800d", x"800d", x"800d", x"800c", x"800c", x"800c", x"800c", 
    x"800c", x"800c", x"800c", x"800c", x"800c", x"800c", x"800c", x"800c", 
    x"800b", x"800b", x"800b", x"800b", x"800b", x"800b", x"800b", x"800b", 
    x"800b", x"800b", x"800b", x"800b", x"800b", x"800a", x"800a", x"800a", 
    x"800a", x"800a", x"800a", x"800a", x"800a", x"800a", x"800a", x"800a", 
    x"800a", x"800a", x"800a", x"8009", x"8009", x"8009", x"8009", x"8009", 
    x"8009", x"8009", x"8009", x"8009", x"8009", x"8009", x"8009", x"8009", 
    x"8009", x"8008", x"8008", x"8008", x"8008", x"8008", x"8008", x"8008", 
    x"8008", x"8008", x"8008", x"8008", x"8008", x"8008", x"8008", x"8008", 
    x"8008", x"8007", x"8007", x"8007", x"8007", x"8007", x"8007", x"8007", 
    x"8007", x"8007", x"8007", x"8007", x"8007", x"8007", x"8007", x"8007", 
    x"8007", x"8006", x"8006", x"8006", x"8006", x"8006", x"8006", x"8006", 
    x"8006", x"8006", x"8006", x"8006", x"8006", x"8006", x"8006", x"8006", 
    x"8006", x"8006", x"8006", x"8006", x"8005", x"8005", x"8005", x"8005", 
    x"8005", x"8005", x"8005", x"8005", x"8005", x"8005", x"8005", x"8005", 
    x"8005", x"8005", x"8005", x"8005", x"8005", x"8005", x"8005", x"8005", 
    x"8004", x"8004", x"8004", x"8004", x"8004", x"8004", x"8004", x"8004", 
    x"8004", x"8004", x"8004", x"8004", x"8004", x"8004", x"8004", x"8004", 
    x"8004", x"8004", x"8004", x"8004", x"8004", x"8004", x"8004", x"8004", 
    x"8003", x"8003", x"8003", x"8003", x"8003", x"8003", x"8003", x"8003", 
    x"8003", x"8003", x"8003", x"8003", x"8003", x"8003", x"8003", x"8003", 
    x"8003", x"8003", x"8003", x"8003", x"8003", x"8003", x"8003", x"8003", 
    x"8003", x"8003", x"8003", x"8003", x"8003", x"8002", x"8002", x"8002", 
    x"8002", x"8002", x"8002", x"8002", x"8002", x"8002", x"8002", x"8002", 
    x"8002", x"8002", x"8002", x"8002", x"8002", x"8002", x"8002", x"8002", 
    x"8002", x"8002", x"8002", x"8002", x"8002", x"8002", x"8002", x"8002", 
    x"8002", x"8002", x"8002", x"8002", x"8002", x"8002", x"8002", x"8002", 
    x"8002", x"8002", x"8002", x"8002", x"8002", x"8002", x"8002", x"8001", 
    x"8001", x"8001", x"8001", x"8001", x"8001", x"8001", x"8001", x"8001", 
    x"8001", x"8001", x"8001", x"8001", x"8001", x"8001", x"8001", x"8001", 
    x"8001", x"8001", x"8001", x"8001", x"8001", x"8001", x"8001", x"8001", 
    x"8001", x"8001", x"8001", x"8001", x"8001", x"8001", x"8001", x"8001", 
    x"8001", x"8001", x"8001", x"8001", x"8001", x"8001", x"8001", x"8001", 
    x"8001", x"8001", x"8001", x"8001", x"8001", x"8001", x"8001", x"8001", 
    x"8001", x"8001", x"8001", x"8001", x"8001", x"8001", x"8001", x"8001");


begin

PROCESS (CLK)
BEGIN
	if (rising_edge (clk)) then
		dADD <= ADD(15);
		msin <= isin(conv_integer(ADD(14 downto 0)));
		mcos <= icos(conv_integer(ADD(14 downto 0)));
		if (dADD = '0') then
			sin <= msin;
			cos <= mcos;
		else
			sin <= x"0" - msin;
			cos <= x"0" - mcos;
		end if;			
	end if;
END PROCESS;


end architecture;
