library IEEE;
use IEEE.std_logic_1164.all; 
use IEEE.std_logic_unsigned.all; 
use ieee.numeric_std.all;

entity bootloader_dp_32 is
  port (
    CLK:              in std_logic;
    WEA:  in std_logic;
    ENA:  in std_logic;
    MASKA:    in std_logic_vector(3 downto 0);
    ADDRA:         in std_logic_vector(11 downto 2);
    DIA:        in std_logic_vector(31 downto 0);
    DOA:         out std_logic_vector(31 downto 0);
    WEB:  in std_logic;
    ENB:  in std_logic;
    ADDRB:         in std_logic_vector(11 downto 2);
    DIB:        in std_logic_vector(31 downto 0);
    MASKB:    in std_logic_vector(3 downto 0);
    DOB:         out std_logic_vector(31 downto 0)
  );
end entity bootloader_dp_32;

architecture behave of bootloader_dp_32 is

  subtype RAM_WORD is STD_LOGIC_VECTOR (31 downto 0);
  type RAM_TABLE is array (0 to 1023) of RAM_WORD;
 shared variable RAM: RAM_TABLE := RAM_TABLE'(
x"0b0b0b99",x"c4040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b99",x"af040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fd0608",x"72830609",x"81058205",x"832b2a83",x"ffff0652",x"04000000",x"00000000",x"00000000",x"71fd0608",x"83ffff73",x"83060981",x"05820583",x"2b2b0906",x"7383ffff",x"0b0b0b0b",x"83a70400",x"72098105",x"72057373",x"09060906",x"73097306",x"070a8106",x"53510400",x"00000000",x"00000000",x"72722473",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71737109",x"71068106",x"30720a10",x"0a720a10",x"0a31050a",x"81065151",x"53510400",x"00000000",x"72722673",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"cc040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"720a722b",x"0a535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72729f06",x"0981050b",x"0b0b88af",x"05040000",x"00000000",x"00000000",x"00000000",x"00000000",x"72722aff",x"739f062a",x"0974090a",x"8106ff05",x"06075351",x"04000000",x"00000000",x"00000000",x"71715351",x"020d0406",x"73830609",x"81058205",x"832b0b2b",x"0772fc06",x"0c515104",x"00000000",x"72098105",x"72050970",x"81050906",x"0a810653",x"51040000",x"00000000",x"00000000",x"00000000",x"72098105",x"72050970",x"81050906",x"0a098106",x"53510400",x"00000000",x"00000000",x"00000000",x"71098105",x"52040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72720981",x"05055351",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097206",x"73730906",x"07535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fc0608",x"72830609",x"81058305",x"1010102a",x"81ff0652",x"04000000",x"00000000",x"00000000",x"71fc0608",x"0b0b0b9c",x"bc738306",x"10100508",x"060b0b0b",x"88b20400",x"00000000",x"00000000",x"0b0b0b89",x"80040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"e8040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097081",x"0509060a",x"8106ff05",x"70547106",x"73097274",x"05ff0506",x"07515151",x"04000000",x"72097081",x"0509060a",x"098106ff",x"05705471",x"06730972",x"7405ff05",x"06075151",x"51040000",x"05ff0504",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"810b0b0b",x"0b9da00c",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71810552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"02840572",x"10100552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"717105ff",x"05715351",x"020d0400",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"81dd3f94",x"8d3f0400",x"00000000",x"00000000",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101053",x"51047381",x"ff067383",x"06098105",x"83051010",x"102b0772",x"fc060c51",x"51043c04",x"72728072",x"8106ff05",x"09720605",x"71105272",x"0a100a53",x"72ed3851",x"51535104",x"88088c08",x"90087575",x"9afd2d50",x"50880856",x"900c8c0c",x"880c5104",x"88088c08",x"90087575",x"9ab92d50",x"50880856",x"900c8c0c",x"880c5104",x"88088c08",x"90088ea6",x"2d900c8c",x"0c880c04",x"ff3d0d0b",x"0b0b9dc4",x"335170a6",x"389dac08",x"70085252",x"70802e92",x"3884129d",x"ac0c702d",x"9dac0870",x"08525270",x"f038810b",x"0b0b0b9d",x"c434833d",x"0d040480",x"3d0d0b0b",x"0b9df008",x"802e8e38",x"0b0b0b0b",x"800b802e",x"09810685",x"38823d0d",x"040b0b0b",x"9df0510b",x"0b0bf5f8",x"3f823d0d",x"0404ff3d",x"0d80c480",x"80845271",x"0870822a",x"70810651",x"515170f3",x"38833d0d",x"04ff3d0d",x"80c48080",x"84527108",x"70812a70",x"81065151",x"5170f338",x"7382900a",x"0c833d0d",x"04fd3d0d",x"75547333",x"7081ff06",x"53537180",x"2e8e3872",x"81ff0651",x"8aa92d81",x"1454e739",x"853d0d04",x"fe3d0d74",x"7080dc80",x"80880c70",x"81ff06ff",x"83115451",x"53718126",x"8d3880fd",x"518aa92d",x"72a03251",x"83397251",x"8aa92d84",x"3d0d0480",x"3d0d83ff",x"ff0b83d0",x"0a0c80fe",x"518aa92d",x"823d0d04",x"ff3d0d83",x"d00a0870",x"882a5252",x"8aec2d71",x"81ff0651",x"8aec2d80",x"fe518aa9",x"2d833d0d",x"0482f6ff",x"0b80cc80",x"80880c80",x"0b80cc80",x"80840c9f",x"0b83900a",x"0c04ff3d",x"0d737008",x"515180c8",x"80808870",x"08708280",x"8007720c",x"5252833d",x"0d04ff3d",x"0d80c880",x"80887008",x"70fdffff",x"06720c52",x"52833d0d",x"04a0900b",x"a0800c9d",x"c80ba084",x"0c99a82d",x"ff3d0d73",x"518b710c",x"90115298",x"8080720c",x"80720c70",x"0883ffff",x"06880c83",x"3d0d04fa",x"3d0d787a",x"7dff1e57",x"57585373",x"ff2ea738",x"80568452",x"75730c72",x"0888180c",x"ff125271",x"f3387484",x"16740872",x"0cff1656",x"565273ff",x"2e098106",x"dd38883d",x"0d04f93d",x"0d80d080",x"80845683",x"d00a0b9c",x"f452588a",x"c92d8c86",x"2d75518c",x"ac2d9dc8",x"70880810",x"10988084",x"05717084",x"05530c56",x"57fb8084",x"a1ad750c",x"9db00b88",x"180c8070",x"770c760c",x"75087083",x"ffff0651",x"5783ffff",x"780ca080",x"54880853",x"77527551",x"8ccb2d75",x"518bea2d",x"77085574",x"772e8938",x"80c3518a",x"a92dff39",x"a0840855",x"74849084",x"b2802e89",x"3880c251",x"8aa92dff",x"399cfc51",x"8ac92d80",x"d00a7008",x"70ffbf06",x"720c5656",x"8a8e2d8c",x"9d2dff3d",x"0d9dd408",x"81119dd4",x"0c518390",x"0a700870",x"feff0672",x"0c525283",x"3d0d0480",x"3d0d8b9b",x"2d728180",x"07518aec",x"2d8bb02d",x"823d0d04",x"fe3d0d80",x"d0808084",x"538c862d",x"85730c80",x"730c7208",x"7081ff06",x"74535152",x"8bea2d71",x"880c843d",x"0d04fc3d",x"0d768111",x"33821233",x"7181800a",x"29718480",x"80290583",x"14337082",x"80291284",x"16335271",x"05a08005",x"86168517",x"33575253",x"53555755",x"53ff1353",x"72ff2e91",x"38737081",x"05553352",x"71757081",x"055734e9",x"3989518e",x"c32d863d",x"0d04f93d",x"0d795780",x"d0808084",x"568c862d",x"81173382",x"18337182",x"80290553",x"5371802e",x"94388517",x"72555372",x"70810554",x"33760cff",x"145473f3",x"38831733",x"84183371",x"82802905",x"56528054",x"73752797",x"38735877",x"760c7317",x"76085353",x"71733481",x"14547474",x"26ed3875",x"518bea2d",x"8b9b2d81",x"84518aec",x"2d74882a",x"518aec2d",x"74518aec",x"2d805473",x"75278f38",x"73177033",x"52528aec",x"2d811454",x"ee398bb0",x"2d893d0d",x"0404fc3d",x"0d768111",x"33821233",x"71902b71",x"882b0783",x"14337072",x"07882b84",x"16337107",x"51525357",x"57545288",x"518ec32d",x"81ff518a",x"a92d80c4",x"80808453",x"72087081",x"2a708106",x"51515271",x"f3387384",x"80800780",x"c4808084",x"0c863d0d",x"04fe3d0d",x"8ed82d88",x"08880881",x"06535371",x"f3388b9b",x"2d818351",x"8aec2d72",x"518aec2d",x"8bb02d84",x"3d0d04fe",x"3d0d800b",x"9dd40c8b",x"9b2d8181",x"518aec2d",x"9db05393",x"52727081",x"05543351",x"8aec2dff",x"125271ff",x"2e098106",x"ec388bb0",x"2d843d0d",x"04fe3d0d",x"800b9dd4",x"0c8b9b2d",x"8182518a",x"ec2d80d0",x"80808453",x"8c862d81",x"d50a0b80",x"d080809c",x"0c80730c",x"72087083",x"b881ff06",x"83b88080",x"07745351",x"528bea2d",x"719ddc0c",x"71902a51",x"8aec2d9d",x"dc08882a",x"518aec2d",x"9ddc0851",x"8aec2d8e",x"d82d8808",x"518aec2d",x"8bb02d84",x"3d0d0480",x"3d0d810b",x"9dd80c80",x"0b83900a",x"0c85518e",x"c32d823d",x"0d04803d",x"0d800b9d",x"d80c8bd1",x"2d86518e",x"c32d823d",x"0d04fd3d",x"0d80d080",x"8084548a",x"518ec32d",x"8c862d9d",x"c8745253",x"8cac2d72",x"88081010",x"98808405",x"71708405",x"530c52fb",x"8084a1ad",x"720c9db0",x"0b88140c",x"73518bea",x"2d8a8e2d",x"8c9d2dfb",x"3d0d80c8",x"8080a852",x"fdffff72",x"08707206",x"740c5253",x"80c88080",x"98700870",x"7506720c",x"52700870",x"fbffff06",x"720c5252",x"f7ffff72",x"08707206",x"740c5272",x"0870efff",x"ff06740c",x"5256dfff",x"ff720870",x"7206740c",x"52720870",x"efff0a06",x"740c5255",x"f7ff0a72",x"08707206",x"740c5272",x"0870fbff",x"0a06740c",x"5254fdff",x"0a720870",x"7206740c",x"525380c8",x"80808870",x"08708480",x"8007720c",x"52700870",x"7806720c",x"52700870",x"90808007",x"720c5270",x"08707706",x"720c5270",x"08709080",x"0a07720c",x"52700870",x"7606720c",x"52700870",x"84800a07",x"720c5270",x"08707506",x"720c5252",x"873d0d04",x"ffab3d0d",x"80d93d08",x"56800b9d",x"d80c800b",x"9dd40c80",x"0bdf8017",x"9db57190",x"2a715656",x"57555772",x"72708105",x"54347388",x"2a537272",x"34738216",x"3475982a",x"52718b16",x"3475902a",x"52718c16",x"3475882a",x"52718d16",x"34758e16",x"348ea60b",x"a0800c80",x"c4808084",x"548480b3",x"740c93e3",x"2d880b80",x"c0808084",x"0c900a53",x"81730c9d",x"94518ac9",x"2d8bd12d",x"fe88880b",x"80dc8080",x"840c81f2",x"0b80d00a",x"0c80d080",x"80847052",x"528bea2d",x"8c862d71",x"518bea2d",x"76777575",x"933d4141",x"5b5b5b83",x"d00a5c78",x"08708106",x"5152719d",x"389dd808",x"5372f038",x"9dd40852",x"87e87227",x"e638727e",x"0c728390",x"0a0c99a1",x"2d82900a",x"08537980",x"2e81b438",x"7280fe2e",x"09810680",x"f4387680",x"2ec13880",x"7d785657",x"5a827727",x"ffb53883",x"ffff7c0c",x"79fe1853",x"53797227",x"983880dc",x"80808872",x"56587216",x"7033790c",x"52811353",x"747326f2",x"38ff1476",x"11547605",x"ff057033",x"74337072",x"882b077f",x"08535155",x"51527173",x"2e098106",x"feed3875",x"3353728a",x"26fee438",x"7210109c",x"c8057652",x"70085152",x"712dfed3",x"397280fd",x"2e098106",x"8638815b",x"fec53976",x"829f269e",x"387a802e",x"87388073",x"a032545b",x"80d73d77",x"05fde005",x"52727234",x"811757fe",x"a239805a",x"fe9d3972",x"80fe2e09",x"8106fe93",x"387957ff",x"7c0c8177",x"5c5afe87",x"398480b3",x"0b80c480",x"80840c04",x"ff3d0d80",x"c4808084",x"52710870",x"812a7081",x"06515151",x"70f33873",x"82900a0c",x"833d0d04",x"ff3d0d80",x"d35198e4",x"2d9a8d2d",x"80cc5198",x"e42d7352",x"805195b0",x"2d833d0d",x"0483fff8",x"0d8d8604",x"83fff80d",x"a0880488",x"0880c080",x"808808a0",x"80082d50",x"880c810b",x"900a0c04",x"98d92dbe",x"0b98e42d",x"5080700c",x"faad95b4",x"da0b8180",x"8071710c",x"7180082e",x"87387011",x"5199d904",x"51bc0b98",x"e42d5099",x"842d0000",x"00000000",x"00000000",x"00000000",x"820b80c0",x"8080900c",x"0b0b0b04",x"0083f00a",x"0b800ba0",x"80721208",x"720c8412",x"5271712e",x"ff05f238",x"028c050d",x"9a800400",x"00000000",x"00000000",x"00000000",x"00fb3d0d",x"77795555",x"80567575",x"24ab3880",x"74249d38",x"80537352",x"745180e1",x"3f880854",x"75802e85",x"38880830",x"5473880c",x"873d0d04",x"73307681",x"325754dc",x"39743055",x"81567380",x"25d238ec",x"39fa3d0d",x"787a5755",x"80577675",x"24a43875",x"9f2c5481",x"53757432",x"74315274",x"519b3f88",x"08547680",x"2e853888",x"08305473",x"880c883d",x"0d047430",x"558157d7",x"39fc3d0d",x"76785354",x"81538074",x"73265255",x"72802e98",x"3870802e",x"a9388072",x"24a43871",x"10731075",x"72265354",x"5272ea38",x"73517883",x"38745170",x"880c863d",x"0d047281",x"2a72812a",x"53537280",x"2ee63871",x"7426ef38",x"73723175",x"74077481",x"2a74812a",x"55555654",x"e539ff3d",x"0d9de40b",x"fc057008",x"525270ff",x"2e913870",x"2dfc1270",x"08525270",x"ff2e0981",x"06f13883",x"3d0d0404",x"ecee3f04",x"00ffffff",x"ff00ffff",x"ffff00ff",x"ffffff00",x"000008df",x"00000911",x"000008b9",x"000007d2",x"00000977",x"0000098e",x"00000865",x"00000866",x"0000077e",x"000009a2",x"43500d0a",x"00000000",x"4c6f6164",x"65642c20",x"73746172",x"74696e67",x"2e2e2e0d",x"0a000000",x"0d0a5a50",x"55494e4f",x"0d0a0000",x"00000000",x"00000000",x"00000000",x"00000eec",x"01090600",x"00000000",x"05b8d800",x"42011900",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"ffffffff",x"00000000",x"ffffffff",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000");

begin

  process (clk)
  begin
    if rising_edge(clk) then
      if ENA='1' then
        if WEA='1' then
          RAM(conv_integer(ADDRA) ) := DIA;
        end if;
        DOA <= RAM(conv_integer(ADDRA)) ;
      end if;
    end if;
  end process;  

  process (clk)
  begin
    if rising_edge(clk) then
      if ENB='1' then
        if WEB='1' then
          RAM( conv_integer(ADDRB) ) := DIB;
        end if;
        DOB <= RAM(conv_integer(ADDRB)) ;
      end if;
    end if;
  end process;  
end behave;
