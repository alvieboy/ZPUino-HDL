library IEEE;
use IEEE.std_logic_1164.all; 
use IEEE.std_logic_unsigned.all; 
use ieee.numeric_std.all;

entity bootloader_dp_32 is
  port (
    CLK:              in std_logic;
    WEA:  in std_logic;
    ENA:  in std_logic;
    MASKA:    in std_logic_vector(3 downto 0);
    ADDRA:         in std_logic_vector(11 downto 2);
    DIA:        in std_logic_vector(31 downto 0);
    DOA:         out std_logic_vector(31 downto 0);
    WEB:  in std_logic;
    ENB:  in std_logic;
    ADDRB:         in std_logic_vector(11 downto 2);
    DIB:        in std_logic_vector(31 downto 0);
    MASKB:    in std_logic_vector(3 downto 0);
    DOB:         out std_logic_vector(31 downto 0)
  );
end entity bootloader_dp_32;

architecture behave of bootloader_dp_32 is

  subtype RAM_WORD is STD_LOGIC_VECTOR (31 downto 0);
  type RAM_TABLE is array (0 to 1023) of RAM_WORD;
 shared variable RAM: RAM_TABLE := RAM_TABLE'(
x"0b0b0b92",x"83040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b89",x"8f040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fd0608",x"72830609",x"81058205",x"832b2a83",x"ffff0652",x"04000000",x"00000000",x"00000000",x"71fd0608",x"83ffff73",x"83060981",x"05820583",x"2b2b0906",x"7383ffff",x"0b0b0b0b",x"83a70400",x"72098105",x"72057373",x"09060906",x"73097306",x"070a8106",x"53510400",x"00000000",x"00000000",x"72722473",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71737109",x"71068106",x"30720a10",x"0a720a10",x"0a31050a",x"81065151",x"53510400",x"00000000",x"72722673",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"c3040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"720a722b",x"0a535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72729f06",x"0981050b",x"0b0b88a6",x"05040000",x"00000000",x"00000000",x"00000000",x"00000000",x"72722aff",x"739f062a",x"0974090a",x"8106ff05",x"06075351",x"04000000",x"00000000",x"00000000",x"71715351",x"020d0406",x"73830609",x"81058205",x"832b0b2b",x"0772fc06",x"0c515104",x"00000000",x"72098105",x"72050970",x"81050906",x"0a810653",x"51040000",x"00000000",x"00000000",x"00000000",x"72098105",x"72050970",x"81050906",x"0a098106",x"53510400",x"00000000",x"00000000",x"00000000",x"71098105",x"52040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72720981",x"05055351",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097206",x"73730906",x"07535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fc0608",x"72830609",x"81058305",x"1010102a",x"81ff0652",x"04000000",x"00000000",x"00000000",x"71fc0608",x"0b0b0b94",x"94738306",x"10100508",x"060b0b0b",x"88a90400",x"00000000",x"00000000",x"0b0b0b88",x"f7040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"df040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097081",x"0509060a",x"8106ff05",x"70547106",x"73097274",x"05ff0506",x"07515151",x"04000000",x"72097081",x"0509060a",x"098106ff",x"05705471",x"06730972",x"7405ff05",x"06075151",x"51040000",x"05ff0504",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"810b0b0b",x"0b97a80c",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71810552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"02840572",x"10100552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"717105ff",x"05715351",x"020d0400",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"81d43f8b",x"e53f0410",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10105351",x"047381ff",x"06738306",x"09810583",x"05101010",x"2b0772fc",x"060c5151",x"043c0472",x"72807281",x"06ff0509",x"72060571",x"1052720a",x"100a5372",x"ed385151",x"53510488",x"088c0890",x"08757592",x"d52d5050",x"88085690",x"0c8c0c88",x"0c510488",x"088c0890",x"08757592",x"912d5050",x"88085690",x"0c8c0c88",x"0c510488",x"088c0890",x"088b9c2d",x"900c8c0c",x"880c04ff",x"3d0d0b0b",x"0b97b833",x"5170a638",x"97b40870",x"08525270",x"802e9238",x"841297b4",x"0c702d97",x"b4087008",x"525270f0",x"38810b0b",x"0b0b97b8",x"34833d0d",x"0404803d",x"0d0b0b0b",x"97d00880",x"2e8e380b",x"0b0b0b80",x"0b802e09",x"81068538",x"823d0d04",x"0b0b0b97",x"d0510b0b",x"0bf6813f",x"823d0d04",x"04ff3d0d",x"80c48080",x"84527108",x"70812a70",x"81065151",x"5170f338",x"7382900a",x"0c833d0d",x"04ff3d0d",x"738f0652",x"89722787",x"3880d712",x"518439b0",x"12518a85",x"2d833d0d",x"04fd3d0d",x"75547333",x"7081ff06",x"53537180",x"2e8e3872",x"81ff0651",x"8a852d81",x"1454e739",x"853d0d04",x"ff3d0d73",x"70842a52",x"528aa52d",x"71518aa5",x"2d833d0d",x"04ff3d0d",x"7370982a",x"52528ae4",x"2d71902a",x"518ae42d",x"71882a51",x"8ae42d71",x"518ae42d",x"833d0d04",x"ff3d0d97",x"bc088111",x"97bc0c51",x"83900a70",x"0870feff",x"06720c52",x"52833d0d",x"04ffb23d",x"0d8480b3",x"0b80c480",x"80840c80",x"c88080a4",x"53fbffff",x"73087072",x"06750c53",x"5480c880",x"80947008",x"70760672",x"0c535380",x"0b80fc80",x"94a45256",x"8ac12d80",x"fc8094c8",x"518ac12d",x"7553fad5",x"aad5aa70",x"740c7308",x"53547174",x"2e098106",x"81f83885",x"aad5aad5",x"70740c73",x"08535471",x"742e0981",x"0681e338",x"faaaeaca",x"da70740c",x"73085354",x"71742e09",x"810681ce",x"3885d7c1",x"d68f7074",x"0c730853",x"5471742e",x"09810681",x"b9388070",x"740c7308",x"53547174",x"2e098106",x"81a838ff",x"70740c73",x"08535471",x"742e0981",x"06819738",x"80d50a70",x"740c7308",x"53547174",x"2e098106",x"81843885",x"a8808070",x"740c7308",x"53547174",x"2e098106",x"80f03882",x"d4807074",x"0c730853",x"5471742e",x"09810680",x"dd3881aa",x"70740c73",x"08535471",x"742e0981",x"0680cb38",x"84135372",x"8880802e",x"098106fe",x"b1387580",x"2e80c038",x"80fc8094",x"e8518ac1",x"2d72518a",x"f92d80fc",x"8094fc51",x"8ac12d73",x"518af92d",x"80fc8095",x"88518ac1",x"2d71518a",x"f92d80fc",x"8094c451",x"8ac12d83",x"f8398156",x"c1398156",x"80ca3980",x"fc809598",x"518ac12d",x"80fc8095",x"b0518ac1",x"2d757654",x"54737370",x"8405550c",x"81145472",x"8880802e",x"098106ed",x"38807055",x"53720852",x"71742e09",x"8106c338",x"81148414",x"54547288",x"80802e09",x"8106e638",x"75802ea0",x"3880fc80",x"94e8518a",x"c12d7251",x"8af92d80",x"fc8094c4",x"518ac12d",x"83873981",x"5680d539",x"80fc8095",x"d0518ac1",x"2d80fc80",x"95f0518a",x"c12d7576",x"56547375",x"70810557",x"34811454",x"74a08080",x"2e098106",x"ed388070",x"55557433",x"7081ff06",x"7581ff06",x"55515271",x"732e0981",x"06ffb838",x"81148116",x"565474a0",x"80802e09",x"8106db38",x"75802ea0",x"3880fc80",x"9698518a",x"c12d7451",x"8af92d80",x"fc8094c4",x"518ac12d",x"828f3981",x"5681c739",x"80fc8096",x"b0518ac1",x"2d80fc80",x"96d0518a",x"c12d7553",x"fad5aad5",x"aa547274",x"740c7308",x"53557174",x"2e098106",x"d23880d5",x"733485ad",x"aad5aa73",x"08535771",x"772e0981",x"06ffbc38",x"81137474",x"0c730853",x"5571742e",x"098106ff",x"aa3880d5",x"7534fad2",x"d6d5aa73",x"08535771",x"772e0981",x"06ff9438",x"81157474",x"0c730853",x"5571742e",x"098106ff",x"823880d5",x"7534fad5",x"a9abaa73",x"08535771",x"772e0981",x"06feec38",x"81157474",x"0c730853",x"5571742e",x"098106fe",x"da3880d5",x"7534fad5",x"aad4d573",x"08535771",x"772e0981",x"06fec438",x"84135372",x"8880802e",x"098106fe",x"d5387580",x"2eb63880",x"fc809698",x"518ac12d",x"74518af9",x"2d80fc80",x"96f4518a",x"c12d7651",x"8af92d80",x"fc809588",x"518ac12d",x"71518af9",x"2d80fc80",x"94c4518a",x"c12d8a39",x"80fc8097",x"84518ac1",x"2dff39ff",x"3d0d8052",x"80518bb9",x"2d833d0d",x"04fb3d0d",x"77795555",x"80567575",x"24ab3880",x"74249d38",x"80537352",x"745180e1",x"3f880854",x"75802e85",x"38880830",x"5473880c",x"873d0d04",x"73307681",x"325754dc",x"39743055",x"81567380",x"25d238ec",x"39fa3d0d",x"787a5755",x"80577675",x"24a43875",x"9f2c5481",x"53757432",x"74315274",x"519b3f88",x"08547680",x"2e853888",x"08305473",x"880c883d",x"0d047430",x"558157d7",x"39fc3d0d",x"76785354",x"81538074",x"73265255",x"72802e98",x"3870802e",x"a9388072",x"24a43871",x"10731075",x"72265354",x"5272ea38",x"73517883",x"38745170",x"880c863d",x"0d047281",x"2a72812a",x"53537280",x"2ee63871",x"7426ef38",x"73723175",x"74077481",x"2a74812a",x"55555654",x"e539ff3d",x"0d97c40b",x"fc057008",x"525270ff",x"2e913870",x"2dfc1270",x"08525270",x"ff2e0981",x"06f13883",x"3d0d0404",x"f58d3f04",x"00ffffff",x"ff00ffff",x"ffff00ff",x"ffffff00",x"5a505569",x"6e6f204d",x"656d6f72",x"79205465",x"73746572",x"20737461",x"7274696e",x"672e0d0a",x"0d0a0000",x"53746172",x"74696e67",x"2073696d",x"706c6520",x"70617474",x"65726e20",x"74657374",x"2e2e2e00",x"4572726f",x"72206174",x"20616464",x"72657373",x"20307800",x"3a207772",x"6f746520",x"30780000",x"2c207265",x"61642062",x"61636b20",x"30780000",x"53746570",x"20312028",x"776f7264",x"29207061",x"73736564",x"2e0d0a00",x"53746172",x"74696e67",x"20696e63",x"72656d65",x"6e74616c",x"20746573",x"742e2e2e",x"00000000",x"53746570",x"20322028",x"696e6372",x"656d656e",x"74616c29",x"20706173",x"7365642e",x"0d0a0000",x"53746172",x"74696e67",x"20627974",x"65776973",x"6520696e",x"6372656d",x"656e7461",x"6c207465",x"73742e2e",x"2e000000",x"0d0a4572",x"726f7220",x"61742061",x"64647265",x"73732030",x"78000000",x"53746570",x"20332028",x"62797465",x"2d776973",x"65292070",x"61737365",x"642e0d0a",x"00000000",x"53746172",x"74696e67",x"20656e64",x"69616e20",x"62797465",x"2d776973",x"65207465",x"73742e2e",x"2e000000",x"3a206578",x"70656374",x"65642030",x"78000000",x"53746570",x"20342028",x"656e6469",x"616e2062",x"7974652d",x"77697365",x"29207061",x"73736564",x"2e0d0a00",x"00000000",x"00000000",x"00000000",x"00000bcc",x"00000000",x"00000000",x"ffffffff",x"00000000",x"ffffffff",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000");

begin

  process (clk)
  begin
    if rising_edge(clk) then
      if ENA='1' then
        if WEA='1' then
          RAM(conv_integer(ADDRA) ) := DIA;
        end if;
        DOA <= RAM(conv_integer(ADDRA)) ;
      end if;
    end if;
  end process;  

  process (clk)
  begin
    if rising_edge(clk) then
      if ENB='1' then
        if WEB='1' then
          RAM( conv_integer(ADDRB) ) := DIB;
        end if;
        DOB <= RAM(conv_integer(ADDRB)) ;
      end if;
    end if;
  end process;  
end behave;
