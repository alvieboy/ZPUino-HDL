--
--  ZPUINO implementation on Spartan3E Evaluation Board from Xilinx
-- 
--  Copyright 2010 Alvaro Lopes <alvieboy@alvie.com>
-- 
--  Version: 1.0
-- 
--  The FreeBSD license
--  
--  Redistribution and use in source and binary forms, with or without
--  modification, are permitted provided that the following conditions
--  are met:
--  
--  1. Redistributions of source code must retain the above copyright
--     notice, this list of conditions and the following disclaimer.
--  2. Redistributions in binary form must reproduce the above
--     copyright notice, this list of conditions and the following
--     disclaimer in the documentation and/or other materials
--     provided with the distribution.
--  
--  THIS SOFTWARE IS PROVIDED BY THE AUTHOR ``AS IS'' AND ANY
--  EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
--  THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
--  PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
--  ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
--  INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
--  (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
--  OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
--  HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
--  STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
--  ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
--  ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
--  
--

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
use work.zpupkg.all;
use work.zpuinopkg.all;
use work.zpuino_config.all;
use work.zpu_config.all;
use work.pad.all;

library UNISIM;
use UNISIM.VCOMPONENTS.all;

entity nexys2_zpuino is
  port (
    CLK         : in    std_logic;
    RST         : in    std_logic;
    UART_RX     : in    std_logic;
    UART_TX     : out   std_logic;
    GPIO        : inout std_logic_vector(zpuino_gpio_count-1 downto 0);
    FPGA_INIT_B : out   std_logic;
    LEDS        : out   std_logic_vector(7 downto 0);

    -- VGA interface
    VGA_RED     : out   std_logic_vector(2 downto 0);
    VGA_GRN     : out   std_logic_vector(2 downto 0);
    VGA_BLU     : out   std_logic_vector(2 downto 1);
    VGA_HS      : out   std_logic;
    VGA_VS      : out   std_logic

  );
end entity nexys2_zpuino;

architecture behave of nexys2_zpuino is

  component clkgen is
  port (
    clkin:  in std_logic;
    rstin:  in std_logic;
    clkout: out std_logic;
    rstout: out std_logic
  );
  end component clkgen;

  component zpuino_serialreset is
  generic (
    SYSTEM_CLOCK_MHZ: integer := 96
  );
  port (
    clk:      in std_logic;
    rx:       in std_logic;
    rstin:    in std_logic;
    rstout:   out std_logic
  );
  end component zpuino_serialreset;



  signal sysrst:      std_logic;
  signal sysclk:      std_logic;
  signal clkgen_rst:  std_logic;

  signal gpio_o: std_logic_vector(zpuino_gpio_count-1 downto 0);
  signal gpio_i: std_logic_vector(zpuino_gpio_count-1 downto 0);
  signal gpio_t: std_logic_vector(zpuino_gpio_count-1 downto 0);

  signal rx: std_logic;
  signal tx: std_logic;

    -- I/O Signals
  signal slot_cyc:   slot_std_logic_type;
  signal slot_we:    slot_std_logic_type;
  signal slot_stb:   slot_std_logic_type;
  signal slot_read:  slot_cpuword_type;
  signal slot_write: slot_cpuword_type;
  signal slot_address:  slot_address_type;
  signal slot_ack:   slot_std_logic_type;
  signal slot_interrupt: slot_std_logic_type;

--  signal spi_enabled:  std_logic;

  signal spi2_enabled:  std_logic;
  signal spi2_mosi:  std_logic;
  signal spi2_miso:  std_logic;
  signal spi2_sck:  std_logic;

--  signal uart_enabled:  std_logic;

  -- SPP signal is one more than GPIO count
  signal gpio_spp_data: std_logic_vector(zpuino_gpio_count-1 downto 0);
  signal gpio_spp_read: std_logic_vector(zpuino_gpio_count-1 downto 0);

  --signal gpio_spp_en: std_logic_vector(zpuino_gpio_count-1 downto 1);

  --signal timers_interrupt:  std_logic_vector(1 downto 0);
  signal timers_spp_data: std_logic_vector(1 downto 0);
  --signal timers_spp_en: std_logic_vector(1 downto 0);
  signal timers_comp: std_logic;

  --signal ivecs: std_logic_vector(17 downto 0);

--  signal sigmadelta_spp_en:  std_logic_vector(1 downto 0);
  signal sigmadelta_spp_data:  std_logic_vector(1 downto 0);

  -- For busy-implementation
--  signal addr_save_q: std_logic_vector(maxAddrBitIncIO downto 0);
  signal write_save_q: std_logic_vector(wordSize-1 downto 0);

  --signal io_address: std_logic_vector(maxAddrBitIncIO downto 0);
  --signal io_write: std_logic_vector(wordSize-1 downto 0);
  --signal io_cyc: std_logic;
  --signal io_stb: std_logic;
  --signal io_we: std_logic;

  --signal io_device_ack: std_logic;

  signal spi_pf_miso: std_logic;
  signal spi_pf_mosi: std_logic;
  signal spi_pf_sck: std_logic;

--  signal adc_mosi:  std_logic;
--  signal adc_miso:  std_logic;
--  signal adc_sck:   std_logic;
-- signal adc_seln:  std_logic;
--  signal adc_enabled: std_logic;

  signal wb_clk_i: std_logic;
  signal wb_rst_i: std_logic;


  -- a 1 in mask bit indicates input capability
  constant spp_cap_in: std_logic_vector(zpuino_gpio_count-1 downto 0) :=
    -- 32 bit word 2 (29 bits used)
    "00000000000000000000000000000" & -- FX2-IO11 - FX2-IO39
    -- 32 bit word 1
    "0000000000" & -- FX2-IO1 - FX2-IO10
    "00" &         -- PS2 CLK/DATA
    "0000" &      -- 4x7-seg LED display, digit anodes, order = AN0-AN3
    "00000000" &  -- 4x7-seg LED display, segment cathodes, order = A,B,C,D,E,F,DP
    "00000000" &  -- Individual LEDs 0-7
    -- 32 bit word 0
    "1" &         -- FX2-IO40
    "000" &       -- pushbuttns BTN1-BTN3
    "1111" &      -- JD dual PMOD connector, pins 1-4 only
    "11111111" &  -- JC dual PMOD connector, pins 1-4, 7-10
    "11111111" &  -- JB dual PMOD connector, pins 1-4, 7-10
    "11111111";   -- JA dual PMOD connector, pins 1-4, 7-10

  -- a 1 in mask bit indicates output capability
  constant spp_cap_out: std_logic_vector(zpuino_gpio_count-1 downto 0) :=
    -- 32 bit word 2 (29 bits used)
    "00000000000000000000000000000" & -- FX2-IO11 - FX2-IO39
    -- 32 bit word 1
    "0000000000" & -- FX2-IO1 - FX2-IO10
    "00" &         -- PS2 CLK/DATA
    "0000" &      -- 4x7-seg LED display, digit anodes, order = AN0-AN3
    "00000000" &  -- 4x7-seg LED display, segment cathodes, order = A,B,C,D,E,F,DP
    "00000000" &  -- Individual LEDs 0-7
    -- 32 bit word 0
    "1" &         -- FX2-IO40
    "000" &       -- pushbuttns BTN1-BTN3
    "1111" &      -- JD dual PMOD connector, pins 1-4 only
    "11111111" &  -- JC dual PMOD connector, pins 1-4, 7-10
    "11111111" &  -- JB dual PMOD connector, pins 1-4, 7-10
    "11111111";   -- JA dual PMOD connector, pins 1-4, 7-10


begin

  wb_clk_i <= sysclk;
  wb_rst_i <= sysrst;

  rstgen: zpuino_serialreset
    generic map (
      SYSTEM_CLOCK_MHZ  => 96
    )
    port map (
      clk       => sysclk,
      rx        => rx,
      rstin     => clkgen_rst,
      rstout    => sysrst
    );

  clkgen_inst: clkgen
  port map (
    clkin   => clk,
    rstin   => rst,
    clkout  => sysclk,
    rstout  => clkgen_rst
  );

  FPGA_INIT_B<='0';


  bufgen:
  for i in 0 to zpuino_gpio_count-1 generate
    iobufgen:
    if spp_cap_out(i) = '1' generate
      iop: IOPAD
        port map(
          I => gpio_o(i),
          O => gpio_i(i),
          T => gpio_t(i),
          C => sysclk,
          PAD => gpio(i)
        );
    end generate iobufgen;
    -- if no output capability, only gen IPAD
    -- to fix bug where GPIO pin is on FPGA input-only pin
    ibufgen:
    if spp_cap_out(i) = '0' generate
      ip: IPAD
        port map(
          O   => gpio_i(i),
          PAD => gpio(i),
          C   => sysclk
        );
    end generate ibufgen;
  end generate;

  ibufrx: IPAD port map ( PAD => UART_RX,  O => rx,  C => sysclk );
  obuftx: OPAD port map ( I => tx,   PAD => UART_TX );

  zpuino:zpuino_top
    port map (
      clk           => sysclk,
      rst           => sysrst,
      slot_cyc      => slot_cyc,
      slot_we       => slot_we,
      slot_stb      => slot_stb,
      slot_read     => slot_read,
      slot_write    => slot_write,
      slot_address  => slot_address,
      slot_ack      => slot_ack,
      slot_interrupt=> slot_interrupt,
      jtag_ctrl_chain_in => (others => '0')
    );

  --
  --
  -- ----------------  I/O connection to devices --------------------
  --
  --

  --
  -- IO SLOT 0
  --

  slot0: zpuino_spi
  port map (
    wb_clk_i  => wb_clk_i,
    wb_rst_i  => wb_rst_i,
    wb_dat_o  => slot_read(0),
    wb_dat_i  => slot_write(0),
    wb_adr_i  => slot_address(0),
    wb_we_i   => slot_we(0),
    wb_cyc_i  => slot_cyc(0),
    wb_stb_i  => slot_stb(0),
    wb_ack_o  => slot_ack(0),
    wb_inta_o => slot_interrupt(0),

    mosi      => spi_pf_mosi,
    miso      => spi_pf_miso,
    sck       => spi_pf_sck,
    enabled   => open--spi_enabled
  );

  --
  -- IO SLOT 1
  --

  uart_inst: zpuino_uart
  port map (
    wb_clk_i  => wb_clk_i,
    wb_rst_i  => wb_rst_i,
    wb_dat_o  => slot_read(1),
    wb_dat_i  => slot_write(1),
    wb_adr_i  => slot_address(1),
    wb_we_i   => slot_we(1),
    wb_cyc_i  => slot_cyc(1),
    wb_stb_i  => slot_stb(1),
    wb_ack_o  => slot_ack(1),

    wb_inta_o => slot_interrupt(1),

    enabled   => open,--uart_enabled,
    tx        => tx,
    rx        => rx
  );

  --
  -- IO SLOT 2
  --

  gpio_inst: zpuino_gpio
  generic map (
    gpio_count => zpuino_gpio_count
  )
  port map (
    wb_clk_i  => wb_clk_i,
    wb_rst_i  => wb_rst_i,
    wb_dat_o  => slot_read(2),
    wb_dat_i  => slot_write(2),
    wb_adr_i  => slot_address(2),
    wb_we_i   => slot_we(2),
    wb_cyc_i  => slot_cyc(2),
    wb_stb_i  => slot_stb(2),
    wb_ack_o  => slot_ack(2),
    wb_inta_o => slot_interrupt(2),

    spp_data  => gpio_spp_data,
    spp_read  => gpio_spp_read,

    gpio_i      => gpio_i,
    gpio_t      => gpio_t,
    gpio_o      => gpio_o,
    spp_cap_in  => spp_cap_in,
    spp_cap_out => spp_cap_out
  );

  --
  -- IO SLOT 3
  --

  timers_inst: zpuino_timers
  port map (
    wb_clk_i  => wb_clk_i,
    wb_rst_i  => wb_rst_i,
    wb_dat_o  => slot_read(3),
    wb_dat_i  => slot_write(3),
    wb_adr_i  => slot_address(3),
    wb_we_i   => slot_we(3),
    wb_cyc_i  => slot_cyc(3),
    wb_stb_i  => slot_stb(3),
    wb_ack_o  => slot_ack(3),

    wb_inta_o => slot_interrupt(3), -- We use two interrupt lines
    wb_intb_o => slot_interrupt(4), -- so we borrow intr line from slot 4

    spp_data  => timers_spp_data,
    spp_en    => open,--timers_spp_en,
    comp      => timers_comp
  );

  --
  -- IO SLOT 4  - DO NOT USE (it's already mapped to Interrupt Controller)
  --

  --
  -- IO SLOT 5
  --

  sigmadelta_inst: zpuino_sigmadelta
  port map (
    wb_clk_i  => wb_clk_i,
    wb_rst_i  => wb_rst_i,
    wb_dat_o  => slot_read(5),
    wb_dat_i  => slot_write(5),
    wb_adr_i  => slot_address(5),
    wb_we_i   => slot_we(5),
    wb_cyc_i  => slot_cyc(5),
    wb_stb_i  => slot_stb(5),
    wb_ack_o  => slot_ack(5),
    wb_inta_o => slot_interrupt(5),

    spp_data  => sigmadelta_spp_data,
    spp_en    => open,--sigmadelta_spp_en,
    sync_in   => timers_comp
  );

  --
  -- IO SLOT 6
  --

  slot1: zpuino_spi
  port map (
    wb_clk_i  => wb_clk_i,
    wb_rst_i  => wb_rst_i,
    wb_dat_o  => slot_read(6),
    wb_dat_i  => slot_write(6),
    wb_adr_i  => slot_address(6),
    wb_we_i   => slot_we(6),
    wb_cyc_i  => slot_cyc(6),
    wb_stb_i  => slot_stb(6),
    wb_ack_o  => slot_ack(6),
    wb_inta_o => slot_interrupt(6),

    mosi      => spi2_mosi,
    miso      => spi2_miso,
    sck       => spi2_sck,
    enabled   => spi2_enabled
  );



  --
  -- IO SLOT 7
  --

  crc16_inst: zpuino_crc16
  port map (
    wb_clk_i  => wb_clk_i,
    wb_rst_i  => wb_rst_i,
    wb_dat_o  => slot_read(7),
    wb_dat_i  => slot_write(7),
    wb_adr_i  => slot_address(7),
    wb_we_i   => slot_we(7),
    wb_cyc_i  => slot_cyc(7),
    wb_stb_i  => slot_stb(7),
    wb_ack_o  => slot_ack(7),
    wb_inta_o => slot_interrupt(7)
  );

  --
  -- IO SLOT 8 (optional)
  --

  adc_inst: zpuino_empty_device
  port map (
    wb_clk_i       => wb_clk_i,
	 	wb_rst_i    => wb_rst_i,
    wb_dat_o      => slot_read(8),
    wb_dat_i     => slot_write(8),
    wb_adr_i   => slot_address(8),
    wb_we_i    => slot_we(8),
    wb_cyc_i      => slot_cyc(8),
    wb_stb_i      => slot_stb(8),
    wb_ack_o      => slot_ack(8),
    wb_inta_o =>  slot_interrupt(8)
  );

  --
  -- IO SLOT 9
  --

  slot9: zpuino_empty_device
  port map (
    wb_clk_i       => wb_clk_i,
	 	wb_rst_i       => wb_rst_i,
    wb_dat_o      => slot_read(9),
    wb_dat_i     => slot_write(9),
    wb_adr_i   => slot_address(9),
    wb_we_i        => slot_we(9),
    wb_cyc_i        => slot_cyc(9),
    wb_stb_i        => slot_stb(9),
    wb_ack_o      => slot_ack(9),
    wb_inta_o => slot_interrupt(9)
  );

  --
  -- IO SLOT 10
  --

  slot10: zpuino_empty_device
  port map (
    wb_clk_i       => wb_clk_i,
	 	wb_rst_i       => wb_rst_i,
    wb_dat_o      => slot_read(10),
    wb_dat_i     => slot_write(10),
    wb_adr_i   => slot_address(10),
    wb_we_i        => slot_we(10),
    wb_cyc_i        => slot_cyc(10),
    wb_stb_i        => slot_stb(10),
    wb_ack_o      => slot_ack(10),
    wb_inta_o => slot_interrupt(10)
  );

  --
  -- IO SLOT 11
  --

  slot11: zpuino_empty_device
  port map (
    wb_clk_i       => wb_clk_i,
	 	wb_rst_i       => wb_rst_i,
    wb_dat_o      => slot_read(11),
    wb_dat_i     => slot_write(11),
    wb_adr_i   => slot_address(11),
    wb_we_i        => slot_we(11),
    wb_cyc_i        => slot_cyc(11),
    wb_stb_i        => slot_stb(11),
    wb_ack_o      => slot_ack(11),
    wb_inta_o => slot_interrupt(11)
  );

  --
  -- IO SLOT 12
  --

  slot12: zpuino_empty_device
  port map (
    wb_clk_i       => wb_clk_i,
	 	wb_rst_i       => wb_rst_i,
    wb_dat_o      => slot_read(12),
    wb_dat_i     => slot_write(12),
    wb_adr_i   => slot_address(12),
    wb_we_i        => slot_we(12),
    wb_cyc_i        => slot_cyc(12),
    wb_stb_i        => slot_stb(12),
    wb_ack_o      => slot_ack(12),
    wb_inta_o => slot_interrupt(12)
  );

  --
  -- IO SLOT 13
  --

  slot13: zpuino_empty_device
  port map (
    wb_clk_i       => wb_clk_i,
	 	wb_rst_i       => wb_rst_i,
    wb_dat_o      => slot_read(13),
    wb_dat_i     => slot_write(13),
    wb_adr_i   => slot_address(13),
    wb_we_i        => slot_we(13),
    wb_cyc_i        => slot_cyc(13),
    wb_stb_i        => slot_stb(13),
    wb_ack_o      => slot_ack(13),
    wb_inta_o => slot_interrupt(13)
  );

  --
  -- IO SLOT 14
  --

  slot14: zpuino_empty_device
  port map (
    wb_clk_i       => wb_clk_i,
	 	wb_rst_i       => wb_rst_i,
    wb_dat_o      => slot_read(14),
    wb_dat_i     => slot_write(14),
    wb_adr_i   => slot_address(14),
    wb_we_i        => slot_we(14),
    wb_cyc_i        => slot_cyc(14),
    wb_stb_i        => slot_stb(14),
    wb_ack_o      => slot_ack(14),
    wb_inta_o => slot_interrupt(14)
  );

  --
  -- IO SLOT 15
  --

  slot15: zpuino_empty_device
  port map (
    wb_clk_i       => wb_clk_i,
	 	wb_rst_i       => wb_rst_i,
    wb_dat_o      => slot_read(15),
    wb_dat_i     => slot_write(15),
    wb_adr_i   => slot_address(15),
    wb_we_i        => slot_we(15),
    wb_cyc_i        => slot_cyc(15),
    wb_stb_i        => slot_stb(15),
    wb_ack_o      => slot_ack(15),
    wb_inta_o => slot_interrupt(15)
  );


  process(
          gpio_spp_read, spi_pf_mosi, spi_pf_sck,
          sigmadelta_spp_data,timers_spp_data,
          spi2_mosi,spi2_sck)
  begin

    gpio_spp_data <= (others => DontCareValue);

    spi_pf_miso <= gpio_spp_read(0);            -- PPS1 : SPI MISO
    gpio_spp_data(1) <= spi_pf_mosi;            -- PPS2 : SPI MOSI
    gpio_spp_data(2) <= spi_pf_sck;             -- PPS3 : SPI SCK
    gpio_spp_data(3) <= sigmadelta_spp_data(0); -- PPS4 : SIGMADELTA DATA
    gpio_spp_data(4) <= timers_spp_data(0);     -- PPS5 : TIMER0
    gpio_spp_data(5) <= timers_spp_data(1);     -- PPS6 : TIMER1
    spi2_miso <= gpio_spp_read(6);              -- PPS7 : USPI MISO
    gpio_spp_data(7) <= spi2_mosi;              -- PPS8 : USPI MOSI
    gpio_spp_data(8) <= spi2_sck;               -- PPS9: USPI SCK
    gpio_spp_data(13) <= sigmadelta_spp_data(1); -- PPS14 : SIGMADELTA1 DATA

    -- External interrupt lines
    --ivecs(16) <= gpio_spp_read(1);
    --ivecs(17) <= gpio_spp_read(2);

  end process;
  
  -- stub off VGA signals for now
  VGA_RED     <= (others => '0');
  VGA_GRN     <= (others => '0');
  VGA_BLU     <= (others => '0');
  VGA_HS      <= '0';
  VGA_VS      <= '0';


end behave;
