library IEEE;
use IEEE.std_logic_1164.all; 
use IEEE.std_logic_unsigned.all; 
use ieee.numeric_std.all;

entity prom_generic_dualport is
  port (
    clk:              in std_logic;
    memAWriteEnable:  in std_logic;
    memAAddr:         in std_logic_vector(14 downto 2);
    memAWrite:        in std_logic_vector(31 downto 0);
    memARead:         out std_logic_vector(31 downto 0);
    memBWriteEnable:  in std_logic;
    memBAddr:         in std_logic_vector(14 downto 2);
    memBWrite:        in std_logic_vector(31 downto 0);
    memBRead:         out std_logic_vector(31 downto 0)
  );
end entity prom_generic_dualport;

architecture behave of prom_generic_dualport is

  subtype RAM_WORD is STD_LOGIC_VECTOR (31 downto 0);
  type RAM_TABLE is array (0 to 8192-1) of RAM_WORD;
  shared variable RAM: RAM_TABLE := RAM_TABLE'(
RAM_WORD'(x"0b0b0ba0"),
RAM_WORD'(x"ac700b0b"),
RAM_WORD'(x"0ba09c0c"),
RAM_WORD'(x"3a0b0b0b"),
RAM_WORD'(x"97840400"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"0b0b0b96"),
RAM_WORD'(x"bf040000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"71fd0608"),
RAM_WORD'(x"72830609"),
RAM_WORD'(x"81058205"),
RAM_WORD'(x"832b2a83"),
RAM_WORD'(x"ffff0652"),
RAM_WORD'(x"04000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"71fd0608"),
RAM_WORD'(x"83ffff73"),
RAM_WORD'(x"83060981"),
RAM_WORD'(x"05820583"),
RAM_WORD'(x"2b2b0906"),
RAM_WORD'(x"7383ffff"),
RAM_WORD'(x"0b0b0b0b"),
RAM_WORD'(x"83a70400"),
RAM_WORD'(x"72098105"),
RAM_WORD'(x"72057373"),
RAM_WORD'(x"09060906"),
RAM_WORD'(x"73097306"),
RAM_WORD'(x"070a8106"),
RAM_WORD'(x"53510400"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"72722473"),
RAM_WORD'(x"732e0753"),
RAM_WORD'(x"51040000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"71737109"),
RAM_WORD'(x"71068106"),
RAM_WORD'(x"30720a10"),
RAM_WORD'(x"0a720a10"),
RAM_WORD'(x"0a31050a"),
RAM_WORD'(x"81065151"),
RAM_WORD'(x"53510400"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"72722673"),
RAM_WORD'(x"732e0753"),
RAM_WORD'(x"51040000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"0b0b0b88"),
RAM_WORD'(x"c3040000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"720a722b"),
RAM_WORD'(x"0a535104"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"72729f06"),
RAM_WORD'(x"0981050b"),
RAM_WORD'(x"0b0b88a6"),
RAM_WORD'(x"05040000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"72722aff"),
RAM_WORD'(x"739f062a"),
RAM_WORD'(x"0974090a"),
RAM_WORD'(x"8106ff05"),
RAM_WORD'(x"06075351"),
RAM_WORD'(x"04000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"71715351"),
RAM_WORD'(x"020d0406"),
RAM_WORD'(x"73830609"),
RAM_WORD'(x"81058205"),
RAM_WORD'(x"832b0b2b"),
RAM_WORD'(x"0772fc06"),
RAM_WORD'(x"0c515104"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"72098105"),
RAM_WORD'(x"72050970"),
RAM_WORD'(x"81050906"),
RAM_WORD'(x"0a810653"),
RAM_WORD'(x"51040000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"72098105"),
RAM_WORD'(x"72050970"),
RAM_WORD'(x"81050906"),
RAM_WORD'(x"0a098106"),
RAM_WORD'(x"53510400"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"71098105"),
RAM_WORD'(x"52040000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"72720981"),
RAM_WORD'(x"05055351"),
RAM_WORD'(x"04000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"72097206"),
RAM_WORD'(x"73730906"),
RAM_WORD'(x"07535104"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"71fc0608"),
RAM_WORD'(x"72830609"),
RAM_WORD'(x"81058305"),
RAM_WORD'(x"1010102a"),
RAM_WORD'(x"81ff0652"),
RAM_WORD'(x"04000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"71fc0608"),
RAM_WORD'(x"0b0b0ba0"),
RAM_WORD'(x"88738306"),
RAM_WORD'(x"10100508"),
RAM_WORD'(x"060b0b0b"),
RAM_WORD'(x"88a90400"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"0b0b0b88"),
RAM_WORD'(x"fe040000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"0b0b0b88"),
RAM_WORD'(x"df040000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"72097081"),
RAM_WORD'(x"0509060a"),
RAM_WORD'(x"8106ff05"),
RAM_WORD'(x"70547106"),
RAM_WORD'(x"73097274"),
RAM_WORD'(x"05ff0506"),
RAM_WORD'(x"07515151"),
RAM_WORD'(x"04000000"),
RAM_WORD'(x"72097081"),
RAM_WORD'(x"0509060a"),
RAM_WORD'(x"098106ff"),
RAM_WORD'(x"05705471"),
RAM_WORD'(x"06730972"),
RAM_WORD'(x"7405ff05"),
RAM_WORD'(x"06075151"),
RAM_WORD'(x"51040000"),
RAM_WORD'(x"05ff0504"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"810b0b0b"),
RAM_WORD'(x"0ba0980c"),
RAM_WORD'(x"51040000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"71810552"),
RAM_WORD'(x"04000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"02840572"),
RAM_WORD'(x"10100552"),
RAM_WORD'(x"04000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"717105ff"),
RAM_WORD'(x"05715351"),
RAM_WORD'(x"020d0400"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"81e83f93"),
RAM_WORD'(x"de3f0410"),
RAM_WORD'(x"10101010"),
RAM_WORD'(x"10101010"),
RAM_WORD'(x"10101010"),
RAM_WORD'(x"10101010"),
RAM_WORD'(x"10101010"),
RAM_WORD'(x"10101010"),
RAM_WORD'(x"10101010"),
RAM_WORD'(x"10105351"),
RAM_WORD'(x"047381ff"),
RAM_WORD'(x"06738306"),
RAM_WORD'(x"09810583"),
RAM_WORD'(x"05101010"),
RAM_WORD'(x"2b0772fc"),
RAM_WORD'(x"060c5151"),
RAM_WORD'(x"043c0472"),
RAM_WORD'(x"72807281"),
RAM_WORD'(x"06ff0509"),
RAM_WORD'(x"72060571"),
RAM_WORD'(x"1052720a"),
RAM_WORD'(x"100a5372"),
RAM_WORD'(x"ed385151"),
RAM_WORD'(x"535104a0"),
RAM_WORD'(x"b008a0b4"),
RAM_WORD'(x"08a0b808"),
RAM_WORD'(x"757598e4"),
RAM_WORD'(x"2d5050a0"),
RAM_WORD'(x"b00856a0"),
RAM_WORD'(x"b80ca0b4"),
RAM_WORD'(x"0ca0b00c"),
RAM_WORD'(x"5104a0b0"),
RAM_WORD'(x"08a0b408"),
RAM_WORD'(x"a0b80875"),
RAM_WORD'(x"7597952d"),
RAM_WORD'(x"5050a0b0"),
RAM_WORD'(x"0856a0b8"),
RAM_WORD'(x"0ca0b40c"),
RAM_WORD'(x"a0b00c51"),
RAM_WORD'(x"04a0b008"),
RAM_WORD'(x"a0b408a0"),
RAM_WORD'(x"b8088bea"),
RAM_WORD'(x"2da0b80c"),
RAM_WORD'(x"a0b40ca0"),
RAM_WORD'(x"b00c04ff"),
RAM_WORD'(x"3d0d0b0b"),
RAM_WORD'(x"0ba0a833"),
RAM_WORD'(x"5170a638"),
RAM_WORD'(x"a0a40870"),
RAM_WORD'(x"08525270"),
RAM_WORD'(x"802e9238"),
RAM_WORD'(x"8412a0a4"),
RAM_WORD'(x"0c702da0"),
RAM_WORD'(x"a4087008"),
RAM_WORD'(x"525270f0"),
RAM_WORD'(x"38810b0b"),
RAM_WORD'(x"0b0ba0a8"),
RAM_WORD'(x"34833d0d"),
RAM_WORD'(x"0404803d"),
RAM_WORD'(x"0d0b0b0b"),
RAM_WORD'(x"9cd80880"),
RAM_WORD'(x"2e8e380b"),
RAM_WORD'(x"0b0b0b80"),
RAM_WORD'(x"0b802e09"),
RAM_WORD'(x"81068538"),
RAM_WORD'(x"823d0d04"),
RAM_WORD'(x"0b0b0b9c"),
RAM_WORD'(x"d8510b0b"),
RAM_WORD'(x"0bf5ed3f"),
RAM_WORD'(x"823d0d04"),
RAM_WORD'(x"04803d0d"),
RAM_WORD'(x"82908408"),
RAM_WORD'(x"70812a70"),
RAM_WORD'(x"81065151"),
RAM_WORD'(x"5170f138"),
RAM_WORD'(x"72829080"),
RAM_WORD'(x"0c823d0d"),
RAM_WORD'(x"04fe3d0d"),
RAM_WORD'(x"747082f0"),
RAM_WORD'(x"880c7081"),
RAM_WORD'(x"ff06ff83"),
RAM_WORD'(x"11545153"),
RAM_WORD'(x"7181268d"),
RAM_WORD'(x"3880fd51"),
RAM_WORD'(x"8a992d72"),
RAM_WORD'(x"a0325183"),
RAM_WORD'(x"3972518a"),
RAM_WORD'(x"992d843d"),
RAM_WORD'(x"0d04ff3d"),
RAM_WORD'(x"0d82f080"),
RAM_WORD'(x"0870882a"),
RAM_WORD'(x"52528ab5"),
RAM_WORD'(x"2d7181ff"),
RAM_WORD'(x"06518ab5"),
RAM_WORD'(x"2d80fe51"),
RAM_WORD'(x"8a992d83"),
RAM_WORD'(x"3d0d0480"),
RAM_WORD'(x"3d0d8290"),
RAM_WORD'(x"840870fb"),
RAM_WORD'(x"ffff0682"),
RAM_WORD'(x"90840c51"),
RAM_WORD'(x"81fff80d"),
RAM_WORD'(x"91be04ff"),
RAM_WORD'(x"39ff3d0d"),
RAM_WORD'(x"82908408"),
RAM_WORD'(x"70810651"),
RAM_WORD'(x"51709f38"),
RAM_WORD'(x"a2f00852"),
RAM_WORD'(x"71ee38a2"),
RAM_WORD'(x"ec085187"),
RAM_WORD'(x"e87127e4"),
RAM_WORD'(x"387182c0"),
RAM_WORD'(x"800c7182"),
RAM_WORD'(x"b0800c8b"),
RAM_WORD'(x"832d8290"),
RAM_WORD'(x"8008a0b0"),
RAM_WORD'(x"0c833d0d"),
RAM_WORD'(x"048386cf"),
RAM_WORD'(x"0b82b088"),
RAM_WORD'(x"0c800b82"),
RAM_WORD'(x"b0840c9f"),
RAM_WORD'(x"0b82b080"),
RAM_WORD'(x"0c04ff3d"),
RAM_WORD'(x"0da2ec08"),
RAM_WORD'(x"8111a2ec"),
RAM_WORD'(x"0c5182b0"),
RAM_WORD'(x"80700870"),
RAM_WORD'(x"feff0672"),
RAM_WORD'(x"0c525283"),
RAM_WORD'(x"3d0d04ff"),
RAM_WORD'(x"3d0d82a0"),
RAM_WORD'(x"84700870"),
RAM_WORD'(x"82800772"),
RAM_WORD'(x"0c525283"),
RAM_WORD'(x"3d0d04ff"),
RAM_WORD'(x"3d0d82a0"),
RAM_WORD'(x"84700870"),
RAM_WORD'(x"fdff0672"),
RAM_WORD'(x"0c525282"),
RAM_WORD'(x"80845185"),
RAM_WORD'(x"710c8071"),
RAM_WORD'(x"0c700870"),
RAM_WORD'(x"81ff0651"),
RAM_WORD'(x"518c872d"),
RAM_WORD'(x"70a0b00c"),
RAM_WORD'(x"833d0d04"),
RAM_WORD'(x"fd3d0d80"),
RAM_WORD'(x"0ba2e808"),
RAM_WORD'(x"53538272"),
RAM_WORD'(x"2784e338"),
RAM_WORD'(x"83ffff0b"),
RAM_WORD'(x"82f0800c"),
RAM_WORD'(x"fe125472"),
RAM_WORD'(x"74278e38"),
RAM_WORD'(x"a0c01333"),
RAM_WORD'(x"82f0880c"),
RAM_WORD'(x"811353ef"),
RAM_WORD'(x"39a2e808"),
RAM_WORD'(x"ff05a2e8"),
RAM_WORD'(x"0ca2e808"),
RAM_WORD'(x"a0c01133"),
RAM_WORD'(x"54ff05a2"),
RAM_WORD'(x"e80ca2e8"),
RAM_WORD'(x"08a0c005"),
RAM_WORD'(x"70337088"),
RAM_WORD'(x"2b750782"),
RAM_WORD'(x"f0800852"),
RAM_WORD'(x"55515271"),
RAM_WORD'(x"732e80cc"),
RAM_WORD'(x"3883ffff"),
RAM_WORD'(x"0b82f080"),
RAM_WORD'(x"0c80fe51"),
RAM_WORD'(x"8a992d81"),
RAM_WORD'(x"ff518ab5"),
RAM_WORD'(x"2d72882a"),
RAM_WORD'(x"518ab52d"),
RAM_WORD'(x"72518ab5"),
RAM_WORD'(x"2d71882a"),
RAM_WORD'(x"518ab52d"),
RAM_WORD'(x"71518ab5"),
RAM_WORD'(x"2d8053a2"),
RAM_WORD'(x"e808732e"),
RAM_WORD'(x"83dd38a0"),
RAM_WORD'(x"c0133351"),
RAM_WORD'(x"8ab52d81"),
RAM_WORD'(x"1353a2e8"),
RAM_WORD'(x"087326ef"),
RAM_WORD'(x"3883c839"),
RAM_WORD'(x"a0c033ff"),
RAM_WORD'(x"05527185"),
RAM_WORD'(x"2683bf38"),
RAM_WORD'(x"7184290b"),
RAM_WORD'(x"0b0b9c90"),
RAM_WORD'(x"05527108"),
RAM_WORD'(x"04800ba2"),
RAM_WORD'(x"ec0c83ff"),
RAM_WORD'(x"ff0b82f0"),
RAM_WORD'(x"800c80fe"),
RAM_WORD'(x"518a992d"),
RAM_WORD'(x"8181518a"),
RAM_WORD'(x"b52d8151"),
RAM_WORD'(x"8ab52d81"),
RAM_WORD'(x"518ab52d"),
RAM_WORD'(x"80518ab5"),
RAM_WORD'(x"2d80518a"),
RAM_WORD'(x"b52d8051"),
RAM_WORD'(x"8ab52d80"),
RAM_WORD'(x"518ab52d"),
RAM_WORD'(x"80ef518a"),
RAM_WORD'(x"b52d81df"),
RAM_WORD'(x"805182e8"),
RAM_WORD'(x"39800ba2"),
RAM_WORD'(x"ec0c83ff"),
RAM_WORD'(x"ff0b82f0"),
RAM_WORD'(x"800c80fe"),
RAM_WORD'(x"518a992d"),
RAM_WORD'(x"8182518a"),
RAM_WORD'(x"b52d82a0"),
RAM_WORD'(x"840870fd"),
RAM_WORD'(x"ff0682a0"),
RAM_WORD'(x"840c5281"),
RAM_WORD'(x"9f0b8280"),
RAM_WORD'(x"840c800b"),
RAM_WORD'(x"8280840c"),
RAM_WORD'(x"800b8280"),
RAM_WORD'(x"840c800b"),
RAM_WORD'(x"8280840c"),
RAM_WORD'(x"82808408"),
RAM_WORD'(x"528c872d"),
RAM_WORD'(x"71902a51"),
RAM_WORD'(x"8ab52d71"),
RAM_WORD'(x"882a518a"),
RAM_WORD'(x"b52d7151"),
RAM_WORD'(x"8ab52d8c"),
RAM_WORD'(x"9b2da0b0"),
RAM_WORD'(x"08518284"),
RAM_WORD'(x"3982a084"),
RAM_WORD'(x"0870fdff"),
RAM_WORD'(x"0682a084"),
RAM_WORD'(x"0c52a0c1"),
RAM_WORD'(x"33a0c233"),
RAM_WORD'(x"71828029"),
RAM_WORD'(x"05535480"),
RAM_WORD'(x"72279638"),
RAM_WORD'(x"a0c57254"),
RAM_WORD'(x"54737081"),
RAM_WORD'(x"05553382"),
RAM_WORD'(x"80840cff"),
RAM_WORD'(x"135372f1"),
RAM_WORD'(x"38a0c333"),
RAM_WORD'(x"a0c43371"),
RAM_WORD'(x"82802905"),
RAM_WORD'(x"55528053"),
RAM_WORD'(x"72742796"),
RAM_WORD'(x"38800b82"),
RAM_WORD'(x"80840c82"),
RAM_WORD'(x"80840852"),
RAM_WORD'(x"71a0c014"),
RAM_WORD'(x"34811353"),
RAM_WORD'(x"e7398c87"),
RAM_WORD'(x"2d83ffff"),
RAM_WORD'(x"0b82f080"),
RAM_WORD'(x"0c80fe51"),
RAM_WORD'(x"8a992d81"),
RAM_WORD'(x"84518ab5"),
RAM_WORD'(x"2d73882a"),
RAM_WORD'(x"518ab52d"),
RAM_WORD'(x"73518ab5"),
RAM_WORD'(x"2d805372"),
RAM_WORD'(x"742780ff"),
RAM_WORD'(x"38a0c013"),
RAM_WORD'(x"33518ab5"),
RAM_WORD'(x"2d811353"),
RAM_WORD'(x"ee39810b"),
RAM_WORD'(x"a2f00c80"),
RAM_WORD'(x"0b82b080"),
RAM_WORD'(x"0c83ffff"),
RAM_WORD'(x"0b82f080"),
RAM_WORD'(x"0c80fe51"),
RAM_WORD'(x"8a992d81"),
RAM_WORD'(x"855180d0"),
RAM_WORD'(x"39800ba2"),
RAM_WORD'(x"f00c8bd5"),
RAM_WORD'(x"2d83ffff"),
RAM_WORD'(x"0b82f080"),
RAM_WORD'(x"0c80fe51"),
RAM_WORD'(x"8a992d81"),
RAM_WORD'(x"8651b539"),
RAM_WORD'(x"82a08408"),
RAM_WORD'(x"70fdff06"),
RAM_WORD'(x"82a0840c"),
RAM_WORD'(x"528c9b2d"),
RAM_WORD'(x"a0b00853"),
RAM_WORD'(x"8c872d72"),
RAM_WORD'(x"81065271"),
RAM_WORD'(x"e33883ff"),
RAM_WORD'(x"ff0b82f0"),
RAM_WORD'(x"800c80fe"),
RAM_WORD'(x"518a992d"),
RAM_WORD'(x"8183518a"),
RAM_WORD'(x"b52d7251"),
RAM_WORD'(x"8ab52d8a"),
RAM_WORD'(x"e22d853d"),
RAM_WORD'(x"0d04fd3d"),
RAM_WORD'(x"0da0800b"),
RAM_WORD'(x"82a08408"),
RAM_WORD'(x"70fdff06"),
RAM_WORD'(x"82a0840c"),
RAM_WORD'(x"52548b0b"),
RAM_WORD'(x"8280840c"),
RAM_WORD'(x"800b8280"),
RAM_WORD'(x"840c800b"),
RAM_WORD'(x"8280840c"),
RAM_WORD'(x"800b8280"),
RAM_WORD'(x"840c800b"),
RAM_WORD'(x"8280840c"),
RAM_WORD'(x"b7df5380"),
RAM_WORD'(x"0b828084"),
RAM_WORD'(x"0c800b82"),
RAM_WORD'(x"80840c80"),
RAM_WORD'(x"0b828084"),
RAM_WORD'(x"0c800b82"),
RAM_WORD'(x"80840c73"),
RAM_WORD'(x"84158280"),
RAM_WORD'(x"8408720c"),
RAM_WORD'(x"ff155555"),
RAM_WORD'(x"5272ff2e"),
RAM_WORD'(x"098106d3"),
RAM_WORD'(x"388c872d"),
RAM_WORD'(x"82808008"),
RAM_WORD'(x"70ffbf06"),
RAM_WORD'(x"8280800c"),
RAM_WORD'(x"5182a080"),
RAM_WORD'(x"0870feff"),
RAM_WORD'(x"0a0682a0"),
RAM_WORD'(x"800c51a0"),
RAM_WORD'(x"880ba080"),
RAM_WORD'(x"0c81fff8"),
RAM_WORD'(x"0da08404"),
RAM_WORD'(x"ff39fd3d"),
RAM_WORD'(x"0d82a090"),
RAM_WORD'(x"53ff730c"),
RAM_WORD'(x"82a09454"),
RAM_WORD'(x"ff740cff"),
RAM_WORD'(x"0b82a098"),
RAM_WORD'(x"0cff0b82"),
RAM_WORD'(x"a09c0c82"),
RAM_WORD'(x"a0847008"),
RAM_WORD'(x"70ef0672"),
RAM_WORD'(x"0c527008"),
RAM_WORD'(x"70a00772"),
RAM_WORD'(x"0c527008"),
RAM_WORD'(x"7080c007"),
RAM_WORD'(x"720c5270"),
RAM_WORD'(x"08708180"),
RAM_WORD'(x"07720c52"),
RAM_WORD'(x"70087082"),
RAM_WORD'(x"8007720c"),
RAM_WORD'(x"5252800b"),
RAM_WORD'(x"82a8800c"),
RAM_WORD'(x"810b82a4"),
RAM_WORD'(x"840c7208"),
RAM_WORD'(x"70fd0674"),
RAM_WORD'(x"0c51830b"),
RAM_WORD'(x"82a48c0c"),
RAM_WORD'(x"720870f7"),
RAM_WORD'(x"06740c51"),
RAM_WORD'(x"840b82a4"),
RAM_WORD'(x"900c7208"),
RAM_WORD'(x"70ef0674"),
RAM_WORD'(x"0c51a80b"),
RAM_WORD'(x"82a5a00c"),
RAM_WORD'(x"730870fd"),
RAM_WORD'(x"ff06750c"),
RAM_WORD'(x"51820b82"),
RAM_WORD'(x"a8880c72"),
RAM_WORD'(x"08708407"),
RAM_WORD'(x"740c51a4"),
RAM_WORD'(x"0b82a590"),
RAM_WORD'(x"0c730870"),
RAM_WORD'(x"ef06750c"),
RAM_WORD'(x"51a50b82"),
RAM_WORD'(x"a5940c73"),
RAM_WORD'(x"0870df06"),
RAM_WORD'(x"750c51a6"),
RAM_WORD'(x"0b82a598"),
RAM_WORD'(x"0c730870"),
RAM_WORD'(x"ffbf0675"),
RAM_WORD'(x"0c51a70b"),
RAM_WORD'(x"82a59c0c"),
RAM_WORD'(x"730870fe"),
RAM_WORD'(x"ff06750c"),
RAM_WORD'(x"51720870"),
RAM_WORD'(x"feff0a06"),
RAM_WORD'(x"740c5182"),
RAM_WORD'(x"a0807008"),
RAM_WORD'(x"7081800a"),
RAM_WORD'(x"07720c52"),
RAM_WORD'(x"730870ff"),
RAM_WORD'(x"bf0a0675"),
RAM_WORD'(x"0c527008"),
RAM_WORD'(x"70ffbf0a"),
RAM_WORD'(x"06720c52"),
RAM_WORD'(x"730870df"),
RAM_WORD'(x"0a06750c"),
RAM_WORD'(x"52700870"),
RAM_WORD'(x"df0a0672"),
RAM_WORD'(x"0c525285"),
RAM_WORD'(x"3d0d04ff"),
RAM_WORD'(x"3d0d800b"),
RAM_WORD'(x"a2f00c80"),
RAM_WORD'(x"0ba2ec0c"),
RAM_WORD'(x"800ba2e8"),
RAM_WORD'(x"0c8bea0b"),
RAM_WORD'(x"a0800c92"),
RAM_WORD'(x"ce2d8481"),
RAM_WORD'(x"d80b8290"),
RAM_WORD'(x"840c810b"),
RAM_WORD'(x"82c0800c"),
RAM_WORD'(x"8bd52d82"),
RAM_WORD'(x"88880b82"),
RAM_WORD'(x"f0840c80"),
RAM_WORD'(x"f20b8280"),
RAM_WORD'(x"800c800b"),
RAM_WORD'(x"a2e40c80"),
RAM_WORD'(x"0ba2e00c"),
RAM_WORD'(x"8b9d2da0"),
RAM_WORD'(x"b008a2e4"),
RAM_WORD'(x"08525270"),
RAM_WORD'(x"802e80e3"),
RAM_WORD'(x"38a0b008"),
RAM_WORD'(x"80fe2e09"),
RAM_WORD'(x"81069238"),
RAM_WORD'(x"a2e80880"),
RAM_WORD'(x"2ede3880"),
RAM_WORD'(x"0ba2e40c"),
RAM_WORD'(x"8cc82dd4"),
RAM_WORD'(x"39a0b008"),
RAM_WORD'(x"80fd2e09"),
RAM_WORD'(x"81068838"),
RAM_WORD'(x"810ba2e0"),
RAM_WORD'(x"0cc239a2"),
RAM_WORD'(x"e8085170"),
RAM_WORD'(x"829f26a3"),
RAM_WORD'(x"38a2e008"),
RAM_WORD'(x"802e8c38"),
RAM_WORD'(x"800ba2e0"),
RAM_WORD'(x"0ca0b008"),
RAM_WORD'(x"a0325271"),
RAM_WORD'(x"a0c01234"),
RAM_WORD'(x"a2e80881"),
RAM_WORD'(x"05a2e80c"),
RAM_WORD'(x"ff963980"),
RAM_WORD'(x"0ba2e40c"),
RAM_WORD'(x"ff8e39a0"),
RAM_WORD'(x"b00880fe"),
RAM_WORD'(x"2e098106"),
RAM_WORD'(x"ff823870"),
RAM_WORD'(x"a2e80c83"),
RAM_WORD'(x"ffff0b82"),
RAM_WORD'(x"f0800c81"),
RAM_WORD'(x"0ba2e40c"),
RAM_WORD'(x"70a2e00c"),
RAM_WORD'(x"feea3980"),
RAM_WORD'(x"3d0da0b0"),
RAM_WORD'(x"08a0b408"),
RAM_WORD'(x"a0b808a0"),
RAM_WORD'(x"80085170"),
RAM_WORD'(x"2da0b80c"),
RAM_WORD'(x"a0b40ca0"),
RAM_WORD'(x"b20c810b"),
RAM_WORD'(x"82c0800c"),
RAM_WORD'(x"823d0d04"),
RAM_WORD'(x"ff3d0d9c"),
RAM_WORD'(x"a80ba088"),
RAM_WORD'(x"52527170"),
RAM_WORD'(x"84055308"),
RAM_WORD'(x"71708405"),
RAM_WORD'(x"530ca0a8"),
RAM_WORD'(x"7126ef38"),
RAM_WORD'(x"833d0d04"),
RAM_WORD'(x"ff3d0d96"),
RAM_WORD'(x"e42d8052"),
RAM_WORD'(x"805194e3"),
RAM_WORD'(x"2d833d0d"),
RAM_WORD'(x"04a0bc08"),
RAM_WORD'(x"02a0bc0c"),
RAM_WORD'(x"f93d0d80"),
RAM_WORD'(x"0ba0bc08"),
RAM_WORD'(x"fc050ca0"),
RAM_WORD'(x"bc088805"),
RAM_WORD'(x"088025b2"),
RAM_WORD'(x"38a0bc08"),
RAM_WORD'(x"88050830"),
RAM_WORD'(x"a0bc0888"),
RAM_WORD'(x"050c800b"),
RAM_WORD'(x"a0bc08f4"),
RAM_WORD'(x"050ca0bc"),
RAM_WORD'(x"08fc0508"),
RAM_WORD'(x"8938810b"),
RAM_WORD'(x"a0bc08f4"),
RAM_WORD'(x"050ca0bc"),
RAM_WORD'(x"08f40508"),
RAM_WORD'(x"a0bc08fc"),
RAM_WORD'(x"050ca0bc"),
RAM_WORD'(x"088c0508"),
RAM_WORD'(x"8025b238"),
RAM_WORD'(x"a0bc088c"),
RAM_WORD'(x"050830a0"),
RAM_WORD'(x"bc088c05"),
RAM_WORD'(x"0c800ba0"),
RAM_WORD'(x"bc08f005"),
RAM_WORD'(x"0ca0bc08"),
RAM_WORD'(x"fc050889"),
RAM_WORD'(x"38810ba0"),
RAM_WORD'(x"bc08f005"),
RAM_WORD'(x"0ca0bc08"),
RAM_WORD'(x"f00508a0"),
RAM_WORD'(x"bc08fc05"),
RAM_WORD'(x"0c8053a0"),
RAM_WORD'(x"bc088c05"),
RAM_WORD'(x"0852a0bc"),
RAM_WORD'(x"08880508"),
RAM_WORD'(x"5181c33f"),
RAM_WORD'(x"a0b00870"),
RAM_WORD'(x"a0bc08f8"),
RAM_WORD'(x"050c54a0"),
RAM_WORD'(x"bc08fc05"),
RAM_WORD'(x"08802e8e"),
RAM_WORD'(x"38a0bc08"),
RAM_WORD'(x"f8050830"),
RAM_WORD'(x"a0bc08f8"),
RAM_WORD'(x"050ca0bc"),
RAM_WORD'(x"08f80508"),
RAM_WORD'(x"70a0b00c"),
RAM_WORD'(x"54893d0d"),
RAM_WORD'(x"a0bc0c04"),
RAM_WORD'(x"a0bc0802"),
RAM_WORD'(x"a0bc0cfb"),
RAM_WORD'(x"3d0d800b"),
RAM_WORD'(x"a0bc08fc"),
RAM_WORD'(x"050ca0bc"),
RAM_WORD'(x"08880508"),
RAM_WORD'(x"80259638"),
RAM_WORD'(x"a0bc0888"),
RAM_WORD'(x"050830a0"),
RAM_WORD'(x"bc088805"),
RAM_WORD'(x"0c810ba0"),
RAM_WORD'(x"bc08fc05"),
RAM_WORD'(x"0ca0bc08"),
RAM_WORD'(x"8c050880"),
RAM_WORD'(x"258e38a0"),
RAM_WORD'(x"bc088c05"),
RAM_WORD'(x"0830a0bc"),
RAM_WORD'(x"088c050c"),
RAM_WORD'(x"8153a0bc"),
RAM_WORD'(x"088c0508"),
RAM_WORD'(x"52a0bc08"),
RAM_WORD'(x"88050851"),
RAM_WORD'(x"b53fa0b0"),
RAM_WORD'(x"0870a0bc"),
RAM_WORD'(x"08f8050c"),
RAM_WORD'(x"54a0bc08"),
RAM_WORD'(x"fc050880"),
RAM_WORD'(x"2e8e38a0"),
RAM_WORD'(x"bc08f805"),
RAM_WORD'(x"0830a0bc"),
RAM_WORD'(x"08f8050c"),
RAM_WORD'(x"a0bc08f8"),
RAM_WORD'(x"050870a0"),
RAM_WORD'(x"b00c5487"),
RAM_WORD'(x"3d0da0bc"),
RAM_WORD'(x"0c04a0bc"),
RAM_WORD'(x"0802a0bc"),
RAM_WORD'(x"0cfd3d0d"),
RAM_WORD'(x"810ba0bc"),
RAM_WORD'(x"08fc050c"),
RAM_WORD'(x"800ba0bc"),
RAM_WORD'(x"08f8050c"),
RAM_WORD'(x"a0bc088c"),
RAM_WORD'(x"0508a0bc"),
RAM_WORD'(x"08880508"),
RAM_WORD'(x"27b238a0"),
RAM_WORD'(x"bc08fc05"),
RAM_WORD'(x"08802ea8"),
RAM_WORD'(x"38800ba0"),
RAM_WORD'(x"bc088c05"),
RAM_WORD'(x"08249d38"),
RAM_WORD'(x"a0bc088c"),
RAM_WORD'(x"050810a0"),
RAM_WORD'(x"bc088c05"),
RAM_WORD'(x"0ca0bc08"),
RAM_WORD'(x"fc050810"),
RAM_WORD'(x"a0bc08fc"),
RAM_WORD'(x"050cc139"),
RAM_WORD'(x"a0bc08fc"),
RAM_WORD'(x"0508802e"),
RAM_WORD'(x"80d538a0"),
RAM_WORD'(x"bc088c05"),
RAM_WORD'(x"08a0bc08"),
RAM_WORD'(x"88050826"),
RAM_WORD'(x"a738a0bc"),
RAM_WORD'(x"08880508"),
RAM_WORD'(x"a0bc088c"),
RAM_WORD'(x"050831a0"),
RAM_WORD'(x"bc088805"),
RAM_WORD'(x"0ca0bc08"),
RAM_WORD'(x"f80508a0"),
RAM_WORD'(x"bc08fc05"),
RAM_WORD'(x"0807a0bc"),
RAM_WORD'(x"08f8050c"),
RAM_WORD'(x"a0bc08fc"),
RAM_WORD'(x"0508812a"),
RAM_WORD'(x"a0bc08fc"),
RAM_WORD'(x"050ca0bc"),
RAM_WORD'(x"088c0508"),
RAM_WORD'(x"812aa0bc"),
RAM_WORD'(x"088c050c"),
RAM_WORD'(x"ffa239a0"),
RAM_WORD'(x"bc089005"),
RAM_WORD'(x"08802e91"),
RAM_WORD'(x"38a0bc08"),
RAM_WORD'(x"88050870"),
RAM_WORD'(x"a0bc08f4"),
RAM_WORD'(x"050c518f"),
RAM_WORD'(x"39a0bc08"),
RAM_WORD'(x"f8050870"),
RAM_WORD'(x"a0bc08f4"),
RAM_WORD'(x"050c51a0"),
RAM_WORD'(x"bc08f405"),
RAM_WORD'(x"08a0b00c"),
RAM_WORD'(x"853d0da0"),
RAM_WORD'(x"bc0c04ff"),
RAM_WORD'(x"3d0d9ccc"),
RAM_WORD'(x"0bfc0570"),
RAM_WORD'(x"08525270"),
RAM_WORD'(x"ff2e9138"),
RAM_WORD'(x"702dfc12"),
RAM_WORD'(x"70085252"),
RAM_WORD'(x"70ff2e09"),
RAM_WORD'(x"8106f138"),
RAM_WORD'(x"833d0d04"),
RAM_WORD'(x"04eda83f"),
RAM_WORD'(x"04000000"),
RAM_WORD'(x"00000709"),
RAM_WORD'(x"0000074d"),
RAM_WORD'(x"00000880"),
RAM_WORD'(x"000007b1"),
RAM_WORD'(x"00000846"),
RAM_WORD'(x"00000865"),
RAM_WORD'(x"00ffffff"),
RAM_WORD'(x"ff00ffff"),
RAM_WORD'(x"ffff00ff"),
RAM_WORD'(x"ffffff00"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000e54"),
RAM_WORD'(x"ffffffff"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"ffffffff"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"0b000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000"),
RAM_WORD'(x"00000000")
);


begin

  process (clk)
  begin
    if rising_edge(clk) then
      if memAWriteEnable='1' then
        RAM( conv_integer(memAAddr) ) := memAWrite;
      end if;
      memARead <= RAM(conv_integer(memAAddr)) ;
    end if;
  end process;  

  process (clk)
  begin
    if rising_edge(clk) then
      if memBWriteEnable='1' then
        RAM( conv_integer(memBAddr) ) := memBWrite;
      end if;
      memBRead <= RAM(conv_integer(memBAddr)) ;
    end if;
  end process;  

end behave; 
