library IEEE;
use IEEE.std_logic_1164.all; 
use IEEE.std_logic_unsigned.all; 
use ieee.numeric_std.all;

entity bootloader_dp_32 is
  port (
    CLK:              in std_logic;
    WEA:  in std_logic;
    ENA:  in std_logic;
    MASKA:    in std_logic_vector(3 downto 0);
    ADDRA:         in std_logic_vector(11 downto 2);
    DIA:        in std_logic_vector(31 downto 0);
    DOA:         out std_logic_vector(31 downto 0);
    WEB:  in std_logic;
    ENB:  in std_logic;
    ADDRB:         in std_logic_vector(11 downto 2);
    DIB:        in std_logic_vector(31 downto 0);
    MASKB:    in std_logic_vector(3 downto 0);
    DOB:         out std_logic_vector(31 downto 0)
  );
end entity bootloader_dp_32;

architecture behave of bootloader_dp_32 is

  subtype RAM_WORD is STD_LOGIC_VECTOR (31 downto 0);
  type RAM_TABLE is array (0 to 1023) of RAM_WORD;
 shared variable RAM: RAM_TABLE := RAM_TABLE'(
x"0b0b0b98",x"c0040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b98",x"a1040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fd0608",x"72830609",x"81058205",x"832b2a83",x"ffff0652",x"04000000",x"00000000",x"00000000",x"71fd0608",x"83ffff73",x"83060981",x"05820583",x"2b2b0906",x"7383ffff",x"0b0b0b0b",x"83a70400",x"72098105",x"72057373",x"09060906",x"73097306",x"070a8106",x"53510400",x"00000000",x"00000000",x"72722473",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71737109",x"71068106",x"30720a10",x"0a720a10",x"0a31050a",x"81065151",x"53510400",x"00000000",x"72722673",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"cc040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"720a722b",x"0a535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72729f06",x"0981050b",x"0b0b88af",x"05040000",x"00000000",x"00000000",x"00000000",x"00000000",x"72722aff",x"739f062a",x"0974090a",x"8106ff05",x"06075351",x"04000000",x"00000000",x"00000000",x"71715351",x"020d0406",x"73830609",x"81058205",x"832b0b2b",x"0772fc06",x"0c515104",x"00000000",x"72098105",x"72050970",x"81050906",x"0a810653",x"51040000",x"00000000",x"00000000",x"00000000",x"72098105",x"72050970",x"81050906",x"0a098106",x"53510400",x"00000000",x"00000000",x"00000000",x"71098105",x"52040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72720981",x"05055351",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097206",x"73730906",x"07535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fc0608",x"72830609",x"81058305",x"1010102a",x"81ff0652",x"04000000",x"00000000",x"00000000",x"71fc0608",x"0b0b0b9e",x"ec738306",x"10100508",x"060b0b0b",x"88b20400",x"00000000",x"00000000",x"0b0b0b89",x"80040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"e8040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097081",x"0509060a",x"8106ff05",x"70547106",x"73097274",x"05ff0506",x"07515151",x"04000000",x"72097081",x"0509060a",x"098106ff",x"05705471",x"06730972",x"7405ff05",x"06075151",x"51040000",x"05ff0504",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"810b0b0b",x"0b9fb40c",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71810552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"02840572",x"10100552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"717105ff",x"05715351",x"020d0400",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"81dd3f96",x"ba3f0400",x"00000000",x"00000000",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101053",x"51047381",x"ff067383",x"06098105",x"83051010",x"102b0772",x"fc060c51",x"51043c04",x"72728072",x"8106ff05",x"09720605",x"71105272",x"0a100a53",x"72ed3851",x"51535104",x"88088c08",x"90087575",x"99ed2d50",x"50880856",x"900c8c0c",x"880c5104",x"88088c08",x"90087575",x"99a92d50",x"50880856",x"900c8c0c",x"880c5104",x"88088c08",x"90088dff",x"2d900c8c",x"0c880c04",x"ff3d0d0b",x"0b0b9fc4",x"335170a6",x"389fc008",x"70085252",x"70802e92",x"3884129f",x"c00c702d",x"9fc00870",x"08525270",x"f038810b",x"0b0b0b9f",x"c434833d",x"0d040480",x"3d0d0b0b",x"0b9ff408",x"802e8e38",x"0b0b0b0b",x"800b802e",x"09810685",x"38823d0d",x"040b0b0b",x"9ff4510b",x"0b0bf5f8",x"3f823d0d",x"0404ff3d",x"0d80c480",x"80845271",x"0870822a",x"70810651",x"515170f3",x"38833d0d",x"04ff3d0d",x"80c48080",x"84527108",x"70812a70",x"81065151",x"5170f338",x"7382900a",x"0c833d0d",x"04fe3d0d",x"747080dc",x"8080880c",x"7081ff06",x"ff831154",x"51537181",x"268d3880",x"fd518aa9",x"2d72a032",x"51833972",x"518aa92d",x"843d0d04",x"803d0d83",x"ffff0b83",x"d00a0c80",x"fe518aa9",x"2d823d0d",x"04ff3d0d",x"83d00a08",x"70882a52",x"528ac92d",x"7181ff06",x"518ac92d",x"80fe518a",x"a92d833d",x"0d0482f6",x"ff0b80cc",x"8080880c",x"800b80cc",x"8080840c",x"9f0b8390",x"0a0c04ff",x"3d0d7370",x"08515180",x"c8808084",x"70087084",x"80800772",x"0c525283",x"3d0d04ff",x"3d0d80c8",x"80808470",x"0870fbff",x"ff06720c",x"5252833d",x"0d04a090",x"0ba0800c",x"9fc80ba0",x"840c98d9",x"2dff3d0d",x"73518b71",x"0c901152",x"98808072",x"0c80720c",x"700883ff",x"ff06880c",x"833d0d04",x"fa3d0d78",x"7a7dff1e",x"57575853",x"73ff2ea7",x"38805684",x"5275730c",x"72088818",x"0cff1252",x"71f33874",x"84167408",x"720cff16",x"56565273",x"ff2e0981",x"06dd3888",x"3d0d04f8",x"3d0d80c0",x"80808457",x"83d00a59",x"8be32d76",x"518c892d",x"9fc87088",x"08101098",x"80840571",x"70840553",x"0c5656fb",x"8084a1ad",x"750c9fa4",x"0b88170c",x"8070780c",x"770c7608",x"83ffff06",x"5683ffdf",x"800b8808",x"278338ff",x"3983ffff",x"790ca080",x"54880853",x"78527651",x"8ca82d76",x"518bc72d",x"78085574",x"762e8938",x"80c3518a",x"a92dff39",x"a0840855",x"74faa090",x"ae802e89",x"3880c251",x"8aa92dff",x"39900a70",x"0870ffbf",x"06720c56",x"568a8e2d",x"8bfa2dff",x"3d0d9fd8",x"0881119f",x"d80c5183",x"900a7008",x"70feff06",x"720c5252",x"833d0d04",x"803d0d8a",x"f82d7281",x"8007518a",x"c92d8b8d",x"2d823d0d",x"04fe3d0d",x"80c08080",x"84538be3",x"2d85730c",x"80730c72",x"087081ff",x"06745351",x"528bc72d",x"71880c84",x"3d0d04fc",x"3d0d7681",x"11338212",x"33718180",x"0a297184",x"80802905",x"83143370",x"82802912",x"84163352",x"7105a080",x"05861685",x"17335752",x"53535557",x"5553ff13",x"5372ff2e",x"91387370",x"81055533",x"52717570",x"81055734",x"e9398951",x"8e9c2d86",x"3d0d04f9",x"3d0d7957",x"80c08080",x"84568be3",x"2d811733",x"82183371",x"82802905",x"53537180",x"2e943885",x"17725553",x"72708105",x"5433760c",x"ff145473",x"f3388317",x"33841833",x"71828029",x"05565280",x"54737527",x"97387358",x"77760c73",x"17760853",x"53717334",x"81145474",x"7426ed38",x"75518bc7",x"2d8af82d",x"8184518a",x"c92d7488",x"2a518ac9",x"2d74518a",x"c92d8054",x"7375278f",x"38731770",x"3352528a",x"c92d8114",x"54ee398b",x"8d2d893d",x"0d04f93d",x"0d795680",x"c0808084",x"558be32d",x"86750c74",x"518bc72d",x"8be32d81",x"ad70760c",x"81173382",x"18337182",x"80290583",x"1933780c",x"84193378",x"0c851933",x"780c5953",x"53805473",x"7727b338",x"72587380",x"2e87388b",x"e32d7775",x"0c731686",x"1133760c",x"87113376",x"0c527451",x"8bc72d8e",x"b12d8808",x"81065271",x"f6388214",x"54767426",x"d1388be3",x"2d84750c",x"74518bc7",x"2d8af82d",x"8187518a",x"c92d8b8d",x"2d893d0d",x"04fc3d0d",x"76811133",x"82123371",x"902b7188",x"2b078314",x"33707207",x"882b8416",x"33710751",x"52535757",x"54528851",x"8e9c2d81",x"ff518aa9",x"2d80c480",x"80845372",x"0870812a",x"70810651",x"515271f3",x"38738480",x"800780c4",x"8080840c",x"863d0d04",x"fe3d0d8e",x"b12d8808",x"88088106",x"535371f3",x"388af82d",x"8183518a",x"c92d7251",x"8ac92d8b",x"8d2d843d",x"0d04fe3d",x"0d800b9f",x"d80c8af8",x"2d818151",x"8ac92d9f",x"a4538f52",x"72708105",x"5433518a",x"c92dff12",x"5271ff2e",x"098106ec",x"388b8d2d",x"843d0d04",x"fe3d0d80",x"0b9fd80c",x"8af82d81",x"82518ac9",x"2d80c080",x"8084528b",x"e32d81f9",x"0a0b80c0",x"80809c0c",x"71087252",x"538bc72d",x"729fe00c",x"72902a51",x"8ac92d9f",x"e008882a",x"518ac92d",x"9fe00851",x"8ac92d8e",x"b12d8808",x"518ac92d",x"8b8d2d84",x"3d0d0480",x"3d0d810b",x"9fdc0c80",x"0b83900a",x"0c85518e",x"9c2d823d",x"0d04803d",x"0d800b9f",x"dc0c8bae",x"2d86518e",x"9c2d823d",x"0d04fd3d",x"0d80c080",x"8084548a",x"518e9c2d",x"8be32d9f",x"c8745253",x"8c892d72",x"88081010",x"98808405",x"71708405",x"530c52fb",x"8084a1ad",x"720c9fa4",x"0b88140c",x"73518bc7",x"2d8a8e2d",x"8bfa2dfc",x"3d0d80c0",x"80808470",x"52558bc7",x"2d8be32d",x"8b750c76",x"80c08080",x"940c8075",x"0ca08054",x"775383d0",x"0a527451",x"8ca82d74",x"518bc72d",x"8a8e2d8b",x"fa2dffab",x"3d0d800b",x"9fdc0c80",x"0b9fd80c",x"800b8dff",x"0ba0800c",x"5780c480",x"80845584",x"80b3750c",x"80c88080",x"a453fbff",x"ff730870",x"7206750c",x"535480c8",x"80809470",x"08707606",x"720c5353",x"a8709aa5",x"71708405",x"530c9b82",x"710c539c",x"9b0b8812",x"0c9daa0b",x"8c120c94",x"bb0b9012",x"0c53880b",x"80d08080",x"840c80d0",x"0a538173",x"0c8bae2d",x"8288880b",x"80dc8080",x"840c81f2",x"0b900a0c",x"80c08080",x"84705252",x"8bc72d8b",x"e32d7151",x"8bc72d8b",x"e32d8472",x"0c71518b",x"c72d7677",x"7675933d",x"41415b5b",x"5b83d00a",x"5c780870",x"81065152",x"719d389f",x"dc085372",x"f0389fd8",x"085287e8",x"7227e638",x"727e0c72",x"83900a0c",x"98d12d82",x"900a0853",x"79802e81",x"b4387280",x"fe2e0981",x"0680f438",x"76802ec1",x"38807d78",x"58565a82",x"7727ffb5",x"3883ffff",x"7c0c79fe",x"18535379",x"72279838",x"80dc8080",x"88725558",x"72157033",x"790c5281",x"13537373",x"26f238ff",x"16751154",x"7505ff05",x"70337433",x"7072882b",x"077f0853",x"51555152",x"71732e09",x"8106feed",x"38743353",x"728a26fe",x"e4387210",x"109ef805",x"75527008",x"5152712d",x"fed33972",x"80fd2e09",x"81068638",x"815bfec5",x"3976829f",x"269e387a",x"802e8738",x"8073a032",x"545b80d7",x"3d7705fd",x"e0055272",x"72348117",x"57fea239",x"805afe9d",x"397280fe",x"2e098106",x"fe933879",x"5783ffff",x"7c0c8177",x"5c5afe85",x"39803d0d",x"88088c08",x"9008a080",x"0851702d",x"900c8c0c",x"8a0c810b",x"80d00a0c",x"823d0d04",x"ff3d0d99",x"882d8052",x"805194f2",x"2d833d0d",x"0483ffff",x"f80d8ce3",x"0483ffff",x"f80d98f0",x"2da08804",x"00000000",x"00000000",x"00000000",x"840b80d0",x"8080900c",x"0b0b0b82",x"0b80d080",x"80900c0b",x"0b0b0400",x"83f00a0b",x"800ba080",x"72120872",x"0c841252",x"71712eff",x"05f23802",x"8c050d98",x"f0040000",x"00fb3d0d",x"77795555",x"80567575",x"24ab3880",x"74249d38",x"80537352",x"745180e1",x"3f880854",x"75802e85",x"38880830",x"5473880c",x"873d0d04",x"73307681",x"325754dc",x"39743055",x"81567380",x"25d238ec",x"39fa3d0d",x"787a5755",x"80577675",x"24a43875",x"9f2c5481",x"53757432",x"74315274",x"519b3f88",x"08547680",x"2e853888",x"08305473",x"880c883d",x"0d047430",x"558157d7",x"39fc3d0d",x"76785354",x"81538074",x"73265255",x"72802e98",x"3870802e",x"a9388072",x"24a43871",x"10731075",x"72265354",x"5272ea38",x"73517883",x"38745170",x"880c863d",x"0d047281",x"2a72812a",x"53537280",x"2ee63871",x"7426ef38",x"73723175",x"74077481",x"2a74812a",x"55555654",x"e539fc3d",x"0d767079",x"7b555555",x"558f7227",x"8c387275",x"07830651",x"70802ea7",x"38ff1252",x"71ff2e98",x"38727081",x"05543374",x"70810556",x"34ff1252",x"71ff2e09",x"8106ea38",x"74880c86",x"3d0d0474",x"51727084",x"05540871",x"70840553",x"0c727084",x"05540871",x"70840553",x"0c727084",x"05540871",x"70840553",x"0c727084",x"05540871",x"70840553",x"0cf01252",x"718f26c9",x"38837227",x"95387270",x"84055408",x"71708405",x"530cfc12",x"52718326",x"ed387054",x"ff8339fc",x"3d0d7679",x"71028c05",x"9f053357",x"55535583",x"72278a38",x"74830651",x"70802ea2",x"38ff1252",x"71ff2e93",x"38737370",x"81055534",x"ff125271",x"ff2e0981",x"06ef3874",x"880c863d",x"0d047474",x"882b7507",x"7071902b",x"07515451",x"8f7227a5",x"38727170",x"8405530c",x"72717084",x"05530c72",x"71708405",x"530c7271",x"70840553",x"0cf01252",x"718f26dd",x"38837227",x"90387271",x"70840553",x"0cfc1252",x"718326f2",x"387053ff",x"9039fb3d",x"0d777970",x"72078306",x"53545270",x"93387173",x"73085456",x"54717308",x"2e80c438",x"73755452",x"71337081",x"ff065254",x"70802e9d",x"38723355",x"70752e09",x"81069538",x"81128114",x"71337081",x"ff065456",x"545270e5",x"38723355",x"7381ff06",x"7581ff06",x"71713188",x"0c525287",x"3d0d0471",x"0970f7fb",x"fdff1406",x"70f88482",x"81800651",x"51517097",x"38841484",x"16710854",x"56547175",x"082edc38",x"73755452",x"ff963980",x"0b880c87",x"3d0d04ff",x"3d0d9fe8",x"0bfc0570",x"08525270",x"ff2e9138",x"702dfc12",x"70085252",x"70ff2e09",x"8106f138",x"833d0d04",x"04eac13f",x"04000000",x"00ffffff",x"ff00ffff",x"ffff00ff",x"ffffff00",x"00000946",x"00000978",x"00000920",x"000007ab",x"000009cf",x"000009e6",x"0000083e",x"000008cd",x"00000757",x"000009fa",x"01090600",x"007fef80",x"05b8d800",x"a4041700",x"00000000",x"00000000",x"00000000",x"00000ff0",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"ffffffff",x"00000000",x"ffffffff",x"00000000",x"00000000",x"00000000",x"00000000");

begin

  process (clk)
  begin
    if rising_edge(clk) then
      if ENA='1' then
        if WEA='1' then
          RAM(conv_integer(ADDRA) ) := DIA;
        end if;
        DOA <= RAM(conv_integer(ADDRA)) ;
      end if;
    end if;
  end process;  

  process (clk)
  begin
    if rising_edge(clk) then
      if ENB='1' then
        if WEB='1' then
          RAM( conv_integer(ADDRB) ) := DIB;
        end if;
        DOB <= RAM(conv_integer(ADDRB)) ;
      end if;
    end if;
  end process;  
end behave;
