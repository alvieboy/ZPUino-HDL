library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;

library work;
use work.zpu_config.all;
use work.zpuino_config.all;
use work.zpupkg.all;
use work.zpuinopkg.all;

library UNISIM;
use UNISIM.vcomponents.all;

entity zpuino_vga_char_ram is
  port (
    -- Scan
    v_clk:    in std_logic;
    v_en:     in std_logic; -- VGA out enable
    v_addr:   in std_logic_vector(11 downto 0); -- Current char
    v_pixel:  out std_logic_vector(7 downto 0); -- Pixel (all 8)

    -- Memory interface
    mi_clk: in std_logic;

    mi_dat_i: in std_logic_vector(7 downto 0); -- Data write
    mi_we:  in std_logic;
    mi_en:  in std_logic;
    mi_dat_o: out std_logic_vector(7 downto 0);
    mi_addr:  in std_logic_vector(11 downto 0)

  );
end entity zpuino_vga_char_ram;


--
--   Address 0 to 15: 1st char
--   Address 16 to 31: 2st char
--
--

architecture behave of zpuino_vga_char_ram is

subtype ramword is std_logic_vector(7 downto 0);

type ramtype is array(0 to 4095) of ramword;

shared variable charram: ramtype := (
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7e",x"81",x"a5",x"81",x"81",x"bd",x"99",x"81",x"81",x"7e",x"00",x"00",x"00",x"00",x"00",x"00",x"7e",x"ff",x"db",x"ff",x"ff",x"c3",x"e7",x"ff",x"ff",x"7e",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6c",x"fe",x"fe",x"fe",x"fe",x"7c",x"38",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"38",x"7c",x"fe",x"7c",x"38",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"3c",x"3c",x"e7",x"e7",x"e7",x"18",x"18",x"3c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"3c",x"7e",x"ff",x"ff",x"7e",x"18",x"18",x"3c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"3c",x"3c",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"e7",x"c3",x"c3",x"e7",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"00",x"00",x"00",x"00",x"00",x"3c",x"66",x"42",x"42",x"66",x"3c",x"00",x"00",x"00",x"00",x"00",x"ff",x"ff",x"ff",x"ff",x"ff",x"c3",x"99",x"bd",x"bd",x"99",x"c3",x"ff",x"ff",x"ff",x"ff",x"ff",x"00",x"00",x"1e",x"0e",x"1a",x"32",x"78",x"cc",x"cc",x"cc",x"cc",x"78",x"00",x"00",x"00",x"00",x"00",x"00",x"3c",x"66",x"66",x"66",x"66",x"3c",x"18",x"7e",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"3f",x"33",x"3f",x"30",x"30",x"30",x"30",x"70",x"f0",x"e0",x"00",x"00",x"00",x"00",x"00",x"00",x"7f",x"63",x"7f",x"63",x"63",x"63",x"63",x"67",x"e7",x"e6",x"c0",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"db",x"3c",x"e7",x"3c",x"db",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"80",x"c0",x"e0",x"f0",x"f8",x"fe",x"f8",x"f0",x"e0",x"c0",x"80",x"00",x"00",x"00",x"00",x"00",x"02",x"06",x"0e",x"1e",x"3e",x"fe",x"3e",x"1e",x"0e",x"06",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"3c",x"7e",x"18",x"18",x"18",x"7e",x"3c",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"00",x"66",x"66",x"00",x"00",x"00",x"00",x"00",x"00",x"7f",x"db",x"db",x"db",x"7b",x"1b",x"1b",x"1b",x"1b",x"1b",x"00",x"00",x"00",x"00",x"00",x"7c",x"c6",x"60",x"38",x"6c",x"c6",x"c6",x"6c",x"38",x"0c",x"c6",x"7c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"fe",x"fe",x"fe",x"fe",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"3c",x"7e",x"18",x"18",x"18",x"7e",x"3c",x"18",x"7e",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"3c",x"7e",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"7e",x"3c",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"0c",x"fe",x"0c",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"30",x"60",x"fe",x"60",x"30",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c0",x"c0",x"c0",x"fe",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"66",x"ff",x"66",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"38",x"38",x"7c",x"7c",x"fe",x"fe",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"fe",x"fe",x"7c",x"7c",x"38",x"38",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"3c",x"3c",x"3c",x"18",x"18",x"18",x"00",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"66",x"66",x"66",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6c",x"6c",x"fe",x"6c",x"6c",x"6c",x"fe",x"6c",x"6c",x"00",x"00",x"00",x"00",x"18",x"18",x"7c",x"c6",x"c2",x"c0",x"7c",x"06",x"06",x"86",x"c6",x"7c",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"c2",x"c6",x"0c",x"18",x"30",x"60",x"c6",x"86",x"00",x"00",x"00",x"00",x"00",x"00",x"38",x"6c",x"6c",x"38",x"76",x"dc",x"cc",x"cc",x"cc",x"76",x"00",x"00",x"00",x"00",x"00",x"30",x"30",x"30",x"60",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0c",x"18",x"30",x"30",x"30",x"30",x"30",x"30",x"18",x"0c",x"00",x"00",x"00",x"00",x"00",x"00",x"30",x"18",x"0c",x"0c",x"0c",x"0c",x"0c",x"0c",x"18",x"30",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"66",x"3c",x"ff",x"3c",x"66",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"7e",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"30",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7e",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"06",x"0c",x"18",x"30",x"60",x"c0",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"7c",x"c6",x"c6",x"ce",x"de",x"f6",x"e6",x"c6",x"c6",x"7c",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"38",x"78",x"18",x"18",x"18",x"18",x"18",x"18",x"7e",x"00",x"00",x"00",x"00",x"00",x"00",x"7c",x"c6",x"06",x"0c",x"18",x"30",x"60",x"c0",x"c6",x"fe",x"00",x"00",x"00",x"00",x"00",x"00",x"7c",x"c6",x"06",x"06",x"3c",x"06",x"06",x"06",x"c6",x"7c",x"00",x"00",x"00",x"00",x"00",x"00",x"0c",x"1c",x"3c",x"6c",x"cc",x"fe",x"0c",x"0c",x"0c",x"1e",x"00",x"00",x"00",x"00",x"00",x"00",x"fe",x"c0",x"c0",x"c0",x"fc",x"06",x"06",x"06",x"c6",x"7c",x"00",x"00",x"00",x"00",x"00",x"00",x"38",x"60",x"c0",x"c0",x"fc",x"c6",x"c6",x"c6",x"c6",x"7c",x"00",x"00",x"00",x"00",x"00",x"00",x"fe",x"c6",x"06",x"06",x"0c",x"18",x"30",x"30",x"30",x"30",x"00",x"00",x"00",x"00",x"00",x"00",x"7c",x"c6",x"c6",x"c6",x"7c",x"c6",x"c6",x"c6",x"c6",x"7c",x"00",x"00",x"00",x"00",x"00",x"00",x"7c",x"c6",x"c6",x"c6",x"7e",x"06",x"06",x"06",x"0c",x"78",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"00",x"00",x"00",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"00",x"00",x"00",x"18",x"18",x"30",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"0c",x"18",x"30",x"60",x"30",x"18",x"0c",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7e",x"00",x"00",x"7e",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"60",x"30",x"18",x"0c",x"06",x"0c",x"18",x"30",x"60",x"00",x"00",x"00",x"00",x"00",x"00",x"7c",x"c6",x"c6",x"0c",x"18",x"18",x"18",x"00",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"7c",x"c6",x"c6",x"c6",x"de",x"de",x"de",x"dc",x"c0",x"7c",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"38",x"6c",x"c6",x"c6",x"fe",x"c6",x"c6",x"c6",x"c6",x"00",x"00",x"00",x"00",x"00",x"00",x"fc",x"66",x"66",x"66",x"7c",x"66",x"66",x"66",x"66",x"fc",x"00",x"00",x"00",x"00",x"00",x"00",x"3c",x"66",x"c2",x"c0",x"c0",x"c0",x"c0",x"c2",x"66",x"3c",x"00",x"00",x"00",x"00",x"00",x"00",x"f8",x"6c",x"66",x"66",x"66",x"66",x"66",x"66",x"6c",x"f8",x"00",x"00",x"00",x"00",x"00",x"00",x"fe",x"66",x"62",x"68",x"78",x"68",x"60",x"62",x"66",x"fe",x"00",x"00",x"00",x"00",x"00",x"00",x"fe",x"66",x"62",x"68",x"78",x"68",x"60",x"60",x"60",x"f0",x"00",x"00",x"00",x"00",x"00",x"00",x"3c",x"66",x"c2",x"c0",x"c0",x"de",x"c6",x"c6",x"66",x"3a",x"00",x"00",x"00",x"00",x"00",x"00",x"c6",x"c6",x"c6",x"c6",x"fe",x"c6",x"c6",x"c6",x"c6",x"c6",x"00",x"00",x"00",x"00",x"00",x"00",x"3c",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"3c",x"00",x"00",x"00",x"00",x"00",x"00",x"1e",x"0c",x"0c",x"0c",x"0c",x"0c",x"cc",x"cc",x"cc",x"78",x"00",x"00",x"00",x"00",x"00",x"00",x"e6",x"66",x"66",x"6c",x"78",x"78",x"6c",x"66",x"66",x"e6",x"00",x"00",x"00",x"00",x"00",x"00",x"f0",x"60",x"60",x"60",x"60",x"60",x"60",x"62",x"66",x"fe",x"00",x"00",x"00",x"00",x"00",x"00",x"c3",x"e7",x"ff",x"ff",x"db",x"c3",x"c3",x"c3",x"c3",x"c3",x"00",x"00",x"00",x"00",x"00",x"00",x"c6",x"e6",x"f6",x"fe",x"de",x"ce",x"c6",x"c6",x"c6",x"c6",x"00",x"00",x"00",x"00",x"00",x"00",x"7c",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"7c",x"00",x"00",x"00",x"00",x"00",x"00",x"fc",x"66",x"66",x"66",x"7c",x"60",x"60",x"60",x"60",x"f0",x"00",x"00",x"00",x"00",x"00",x"00",x"7c",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"d6",x"de",x"7c",x"0c",x"0e",x"00",x"00",x"00",x"00",x"fc",x"66",x"66",x"66",x"7c",x"6c",x"66",x"66",x"66",x"e6",x"00",x"00",x"00",x"00",x"00",x"00",x"7c",x"c6",x"c6",x"60",x"38",x"0c",x"06",x"c6",x"c6",x"7c",x"00",x"00",x"00",x"00",x"00",x"00",x"ff",x"db",x"99",x"18",x"18",x"18",x"18",x"18",x"18",x"3c",x"00",x"00",x"00",x"00",x"00",x"00",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"7c",x"00",x"00",x"00",x"00",x"00",x"00",x"c3",x"c3",x"c3",x"c3",x"c3",x"c3",x"c3",x"66",x"3c",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"c3",x"c3",x"c3",x"c3",x"c3",x"db",x"db",x"ff",x"66",x"66",x"00",x"00",x"00",x"00",x"00",x"00",x"c3",x"c3",x"66",x"3c",x"18",x"18",x"3c",x"66",x"c3",x"c3",x"00",x"00",x"00",x"00",x"00",x"00",x"c3",x"c3",x"c3",x"66",x"3c",x"18",x"18",x"18",x"18",x"3c",x"00",x"00",x"00",x"00",x"00",x"00",x"ff",x"c3",x"86",x"0c",x"18",x"30",x"60",x"c1",x"c3",x"ff",x"00",x"00",x"00",x"00",x"00",x"00",x"3c",x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"3c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"c0",x"e0",x"70",x"38",x"1c",x"0e",x"06",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"3c",x"0c",x"0c",x"0c",x"0c",x"0c",x"0c",x"0c",x"0c",x"3c",x"00",x"00",x"00",x"00",x"10",x"38",x"6c",x"c6",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"ff",x"00",x"00",x"30",x"30",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"78",x"0c",x"7c",x"cc",x"cc",x"cc",x"76",x"00",x"00",x"00",x"00",x"00",x"00",x"e0",x"60",x"60",x"78",x"6c",x"66",x"66",x"66",x"66",x"7c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7c",x"c6",x"c0",x"c0",x"c0",x"c6",x"7c",x"00",x"00",x"00",x"00",x"00",x"00",x"1c",x"0c",x"0c",x"3c",x"6c",x"cc",x"cc",x"cc",x"cc",x"76",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7c",x"c6",x"fe",x"c0",x"c0",x"c6",x"7c",x"00",x"00",x"00",x"00",x"00",x"00",x"38",x"6c",x"64",x"60",x"f0",x"60",x"60",x"60",x"60",x"f0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"76",x"cc",x"cc",x"cc",x"cc",x"cc",x"7c",x"0c",x"cc",x"78",x"00",x"00",x"00",x"e0",x"60",x"60",x"6c",x"76",x"66",x"66",x"66",x"66",x"e6",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"00",x"38",x"18",x"18",x"18",x"18",x"18",x"3c",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"06",x"00",x"0e",x"06",x"06",x"06",x"06",x"06",x"06",x"66",x"66",x"3c",x"00",x"00",x"00",x"e0",x"60",x"60",x"66",x"6c",x"78",x"78",x"6c",x"66",x"e6",x"00",x"00",x"00",x"00",x"00",x"00",x"38",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"3c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"e6",x"ff",x"db",x"db",x"db",x"db",x"db",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"dc",x"66",x"66",x"66",x"66",x"66",x"66",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7c",x"c6",x"c6",x"c6",x"c6",x"c6",x"7c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"dc",x"66",x"66",x"66",x"66",x"66",x"7c",x"60",x"60",x"f0",x"00",x"00",x"00",x"00",x"00",x"00",x"76",x"cc",x"cc",x"cc",x"cc",x"cc",x"7c",x"0c",x"0c",x"1e",x"00",x"00",x"00",x"00",x"00",x"00",x"dc",x"76",x"66",x"60",x"60",x"60",x"f0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7c",x"c6",x"60",x"38",x"0c",x"c6",x"7c",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"30",x"30",x"fc",x"30",x"30",x"30",x"30",x"36",x"1c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"76",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c3",x"c3",x"c3",x"c3",x"66",x"3c",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c3",x"c3",x"c3",x"db",x"db",x"ff",x"66",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c3",x"66",x"3c",x"18",x"3c",x"66",x"c3",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"7e",x"06",x"0c",x"f8",x"00",x"00",x"00",x"00",x"00",x"00",x"fe",x"cc",x"18",x"30",x"60",x"c6",x"fe",x"00",x"00",x"00",x"00",x"00",x"00",x"0e",x"18",x"18",x"18",x"70",x"18",x"18",x"18",x"18",x"0e",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"00",x"18",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"70",x"18",x"18",x"18",x"0e",x"18",x"18",x"18",x"18",x"70",x"00",x"00",x"00",x"00",x"00",x"00",x"76",x"dc",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"38",x"6c",x"c6",x"c6",x"c6",x"fe",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3c",x"66",x"c2",x"c0",x"c0",x"c0",x"c2",x"66",x"3c",x"0c",x"06",x"7c",x"00",x"00",x"00",x"00",x"cc",x"00",x"00",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"76",x"00",x"00",x"00",x"00",x"00",x"0c",x"18",x"30",x"00",x"7c",x"c6",x"fe",x"c0",x"c0",x"c6",x"7c",x"00",x"00",x"00",x"00",x"00",x"10",x"38",x"6c",x"00",x"78",x"0c",x"7c",x"cc",x"cc",x"cc",x"76",x"00",x"00",x"00",x"00",x"00",x"00",x"cc",x"00",x"00",x"78",x"0c",x"7c",x"cc",x"cc",x"cc",x"76",x"00",x"00",x"00",x"00",x"00",x"60",x"30",x"18",x"00",x"78",x"0c",x"7c",x"cc",x"cc",x"cc",x"76",x"00",x"00",x"00",x"00",x"00",x"38",x"6c",x"38",x"00",x"78",x"0c",x"7c",x"cc",x"cc",x"cc",x"76",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3c",x"66",x"60",x"60",x"66",x"3c",x"0c",x"06",x"3c",x"00",x"00",x"00",x"00",x"10",x"38",x"6c",x"00",x"7c",x"c6",x"fe",x"c0",x"c0",x"c6",x"7c",x"00",x"00",x"00",x"00",x"00",x"00",x"c6",x"00",x"00",x"7c",x"c6",x"fe",x"c0",x"c0",x"c6",x"7c",x"00",x"00",x"00",x"00",x"00",x"60",x"30",x"18",x"00",x"7c",x"c6",x"fe",x"c0",x"c0",x"c6",x"7c",x"00",x"00",x"00",x"00",x"00",x"00",x"66",x"00",x"00",x"38",x"18",x"18",x"18",x"18",x"18",x"3c",x"00",x"00",x"00",x"00",x"00",x"18",x"3c",x"66",x"00",x"38",x"18",x"18",x"18",x"18",x"18",x"3c",x"00",x"00",x"00",x"00",x"00",x"60",x"30",x"18",x"00",x"38",x"18",x"18",x"18",x"18",x"18",x"3c",x"00",x"00",x"00",x"00",x"00",x"c6",x"00",x"10",x"38",x"6c",x"c6",x"c6",x"fe",x"c6",x"c6",x"c6",x"00",x"00",x"00",x"00",x"38",x"6c",x"38",x"00",x"38",x"6c",x"c6",x"c6",x"fe",x"c6",x"c6",x"c6",x"00",x"00",x"00",x"00",x"18",x"30",x"60",x"00",x"fe",x"66",x"60",x"7c",x"60",x"60",x"66",x"fe",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6e",x"3b",x"1b",x"7e",x"d8",x"dc",x"77",x"00",x"00",x"00",x"00",x"00",x"00",x"3e",x"6c",x"cc",x"cc",x"fe",x"cc",x"cc",x"cc",x"cc",x"ce",x"00",x"00",x"00",x"00",x"00",x"10",x"38",x"6c",x"00",x"7c",x"c6",x"c6",x"c6",x"c6",x"c6",x"7c",x"00",x"00",x"00",x"00",x"00",x"00",x"c6",x"00",x"00",x"7c",x"c6",x"c6",x"c6",x"c6",x"c6",x"7c",x"00",x"00",x"00",x"00",x"00",x"60",x"30",x"18",x"00",x"7c",x"c6",x"c6",x"c6",x"c6",x"c6",x"7c",x"00",x"00",x"00",x"00",x"00",x"30",x"78",x"cc",x"00",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"76",x"00",x"00",x"00",x"00",x"00",x"60",x"30",x"18",x"00",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"76",x"00",x"00",x"00",x"00",x"00",x"00",x"c6",x"00",x"00",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"7e",x"06",x"0c",x"78",x"00",x"00",x"c6",x"00",x"7c",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"7c",x"00",x"00",x"00",x"00",x"00",x"c6",x"00",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"7c",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"7e",x"c3",x"c0",x"c0",x"c0",x"c3",x"7e",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"38",x"6c",x"64",x"60",x"f0",x"60",x"60",x"60",x"60",x"e6",x"fc",x"00",x"00",x"00",x"00",x"00",x"00",x"c3",x"66",x"3c",x"18",x"ff",x"18",x"ff",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"fc",x"66",x"66",x"7c",x"62",x"66",x"6f",x"66",x"66",x"66",x"f3",x"00",x"00",x"00",x"00",x"00",x"0e",x"1b",x"18",x"18",x"18",x"7e",x"18",x"18",x"18",x"18",x"18",x"d8",x"70",x"00",x"00",x"00",x"18",x"30",x"60",x"00",x"78",x"0c",x"7c",x"cc",x"cc",x"cc",x"76",x"00",x"00",x"00",x"00",x"00",x"0c",x"18",x"30",x"00",x"38",x"18",x"18",x"18",x"18",x"18",x"3c",x"00",x"00",x"00",x"00",x"00",x"18",x"30",x"60",x"00",x"7c",x"c6",x"c6",x"c6",x"c6",x"c6",x"7c",x"00",x"00",x"00",x"00",x"00",x"18",x"30",x"60",x"00",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"76",x"00",x"00",x"00",x"00",x"00",x"00",x"76",x"dc",x"00",x"dc",x"66",x"66",x"66",x"66",x"66",x"66",x"00",x"00",x"00",x"00",x"76",x"dc",x"00",x"c6",x"e6",x"f6",x"fe",x"de",x"ce",x"c6",x"c6",x"c6",x"00",x"00",x"00",x"00",x"00",x"3c",x"6c",x"6c",x"3e",x"00",x"7e",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"38",x"6c",x"6c",x"38",x"00",x"7c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"30",x"30",x"00",x"30",x"30",x"60",x"c0",x"c6",x"c6",x"7c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"fe",x"c0",x"c0",x"c0",x"c0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"fe",x"06",x"06",x"06",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"c0",x"c0",x"c2",x"c6",x"cc",x"18",x"30",x"60",x"ce",x"9b",x"06",x"0c",x"1f",x"00",x"00",x"00",x"c0",x"c0",x"c2",x"c6",x"cc",x"18",x"30",x"66",x"ce",x"96",x"3e",x"06",x"06",x"00",x"00",x"00",x"00",x"18",x"18",x"00",x"18",x"18",x"18",x"3c",x"3c",x"3c",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"36",x"6c",x"d8",x"6c",x"36",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"d8",x"6c",x"36",x"6c",x"d8",x"00",x"00",x"00",x"00",x"00",x"00",x"11",x"44",x"11",x"44",x"11",x"44",x"11",x"44",x"11",x"44",x"11",x"44",x"11",x"44",x"11",x"44",x"55",x"aa",x"55",x"aa",x"55",x"aa",x"55",x"aa",x"55",x"aa",x"55",x"aa",x"55",x"aa",x"55",x"aa",x"dd",x"77",x"dd",x"77",x"dd",x"77",x"dd",x"77",x"dd",x"77",x"dd",x"77",x"dd",x"77",x"dd",x"77",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"f8",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"f8",x"18",x"f8",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"f6",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"fe",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"00",x"00",x"00",x"00",x"00",x"f8",x"18",x"f8",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"36",x"36",x"36",x"36",x"36",x"f6",x"06",x"f6",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"00",x"00",x"00",x"00",x"00",x"fe",x"06",x"f6",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"f6",x"06",x"fe",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"fe",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"18",x"f8",x"18",x"f8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"f8",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"1f",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"ff",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"ff",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"1f",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"ff",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"ff",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"1f",x"18",x"1f",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"37",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"37",x"30",x"3f",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3f",x"30",x"37",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"f7",x"00",x"ff",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"ff",x"00",x"f7",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"37",x"30",x"37",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"00",x"00",x"00",x"00",x"00",x"ff",x"00",x"ff",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"36",x"36",x"36",x"36",x"36",x"f7",x"00",x"f7",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"18",x"18",x"18",x"18",x"18",x"ff",x"00",x"ff",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"ff",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"ff",x"00",x"ff",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"ff",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"3f",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"18",x"1f",x"18",x"1f",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"1f",x"18",x"1f",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3f",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"ff",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"18",x"18",x"18",x"18",x"18",x"ff",x"18",x"ff",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"f8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"1f",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"0f",x"0f",x"0f",x"0f",x"0f",x"0f",x"0f",x"0f",x"0f",x"0f",x"0f",x"0f",x"0f",x"0f",x"0f",x"0f",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"76",x"dc",x"d8",x"d8",x"d8",x"dc",x"76",x"00",x"00",x"00",x"00",x"00",x"00",x"78",x"cc",x"cc",x"cc",x"d8",x"cc",x"c6",x"c6",x"c6",x"cc",x"00",x"00",x"00",x"00",x"00",x"00",x"fe",x"c6",x"c6",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"fe",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"fe",x"c6",x"60",x"30",x"18",x"30",x"60",x"c6",x"fe",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7e",x"d8",x"d8",x"d8",x"d8",x"d8",x"70",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"66",x"66",x"66",x"66",x"66",x"7c",x"60",x"60",x"c0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"76",x"dc",x"18",x"18",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7e",x"18",x"3c",x"66",x"66",x"66",x"3c",x"18",x"7e",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"38",x"6c",x"c6",x"c6",x"fe",x"c6",x"c6",x"6c",x"38",x"00",x"00",x"00",x"00",x"00",x"00",x"38",x"6c",x"c6",x"c6",x"c6",x"6c",x"6c",x"6c",x"6c",x"ee",x"00",x"00",x"00",x"00",x"00",x"00",x"1e",x"30",x"18",x"0c",x"3e",x"66",x"66",x"66",x"66",x"3c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7e",x"db",x"db",x"db",x"7e",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"06",x"7e",x"db",x"db",x"f3",x"7e",x"60",x"c0",x"00",x"00",x"00",x"00",x"00",x"00",x"1c",x"30",x"60",x"60",x"7c",x"60",x"60",x"60",x"30",x"1c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7c",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"fe",x"00",x"00",x"fe",x"00",x"00",x"fe",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"7e",x"18",x"18",x"00",x"00",x"ff",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"30",x"18",x"0c",x"06",x"0c",x"18",x"30",x"00",x"7e",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0c",x"18",x"30",x"60",x"30",x"18",x"0c",x"00",x"7e",x"00",x"00",x"00",x"00",x"00",x"00",x"0e",x"1b",x"1b",x"1b",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"d8",x"d8",x"d8",x"70",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"00",x"7e",x"00",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"76",x"dc",x"00",x"76",x"dc",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"38",x"6c",x"6c",x"38",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0f",x"0c",x"0c",x"0c",x"0c",x"0c",x"ec",x"6c",x"6c",x"3c",x"1c",x"00",x"00",x"00",x"00",x"00",x"d8",x"6c",x"6c",x"6c",x"6c",x"6c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"70",x"d8",x"30",x"60",x"c8",x"f8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7c",x"7c",x"7c",x"7c",x"7c",x"7c",x"7c",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
);

begin

  -- VGA port
  process(v_clk)
  begin
    if rising_edge(v_clk) then
      if v_en='1' then
        v_pixel <= charram(conv_integer(v_addr));
      end if;
    end if;
  end process;

  
  -- CPU interface
  process(mi_clk)
  begin
    if rising_edge(mi_clk) then
      if mi_en='1' then
        if mi_we='1' then
          charram(conv_integer(mi_addr)):=mi_dat_i;
        end if;
        mi_dat_o <= charram(conv_integer(mi_addr));
      end if;
    end if;
  end process;

end behave;
