library IEEE;
use IEEE.std_logic_1164.all; 
use IEEE.std_logic_unsigned.all; 
use ieee.numeric_std.all;

entity bootloader_dp_32 is
  port (
    CLK:              in std_logic;
    WEA:  in std_logic;
    ENA:  in std_logic;
    MASKA:    in std_logic_vector(3 downto 0);
    ADDRA:         in std_logic_vector(11 downto 2);
    DIA:        in std_logic_vector(31 downto 0);
    DOA:         out std_logic_vector(31 downto 0);
    WEB:  in std_logic;
    ENB:  in std_logic;
    ADDRB:         in std_logic_vector(11 downto 2);
    DIB:        in std_logic_vector(31 downto 0);
    MASKB:    in std_logic_vector(3 downto 0);
    DOB:         out std_logic_vector(31 downto 0)
  );
end entity bootloader_dp_32;

architecture behave of bootloader_dp_32 is

  subtype RAM_WORD is STD_LOGIC_VECTOR (31 downto 0);
  type RAM_TABLE is array (0 to 1023) of RAM_WORD;
 shared variable RAM: RAM_TABLE := RAM_TABLE'(
x"0b0b0b9b",x"b5040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b9b",x"a0040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fd0608",x"72830609",x"81058205",x"832b2a83",x"ffff0652",x"04000000",x"00000000",x"00000000",x"71fd0608",x"83ffff73",x"83060981",x"05820583",x"2b2b0906",x"7383ffff",x"0b0b0b0b",x"83a70400",x"72098105",x"72057373",x"09060906",x"73097306",x"070a8106",x"53510400",x"00000000",x"00000000",x"72722473",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71737109",x"71068106",x"30720a10",x"0a720a10",x"0a31050a",x"81065151",x"53510400",x"00000000",x"72722673",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"cc040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"720a722b",x"0a535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72729f06",x"0981050b",x"0b0b88af",x"05040000",x"00000000",x"00000000",x"00000000",x"00000000",x"72722aff",x"739f062a",x"0974090a",x"8106ff05",x"06075351",x"04000000",x"00000000",x"00000000",x"71715351",x"020d0406",x"73830609",x"81058205",x"832b0b2b",x"0772fc06",x"0c515104",x"00000000",x"72098105",x"72050970",x"81050906",x"0a810653",x"51040000",x"00000000",x"00000000",x"00000000",x"72098105",x"72050970",x"81050906",x"0a098106",x"53510400",x"00000000",x"00000000",x"00000000",x"71098105",x"52040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72720981",x"05055351",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097206",x"73730906",x"07535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fc0608",x"72830609",x"81058305",x"1010102a",x"81ff0652",x"04000000",x"00000000",x"00000000",x"71fc0608",x"0b0b0b9d",x"fc738306",x"10100508",x"060b0b0b",x"88b20400",x"00000000",x"00000000",x"0b0b0b89",x"80040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"e8040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097081",x"0509060a",x"8106ff05",x"70547106",x"73097274",x"05ff0506",x"07515151",x"04000000",x"72097081",x"0509060a",x"098106ff",x"05705471",x"06730972",x"7405ff05",x"06075151",x"51040000",x"05ff0504",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"810b0b0b",x"0b9ec00c",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71810552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"02840572",x"10100552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"717105ff",x"05715351",x"020d0400",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"81d53f95",x"d53f0400",x"00000000",x"00000000",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101053",x"51047381",x"ff067383",x"06098105",x"83051010",x"102b0772",x"fc060c51",x"51043c04",x"72728072",x"8106ff05",x"09720605",x"71105272",x"0a100a53",x"72ed3851",x"51535104",x"88088c08",x"90087575",x"9cd42d50",x"50880856",x"900c8c0c",x"880c5104",x"88088c08",x"90087575",x"9c992d50",x"50880856",x"900c8c0c",x"880c5104",x"88088c08",x"90088eb1",x"2d900c8c",x"0c880c04",x"ff3d0d0b",x"0b0b9ee4",x"3351709e",x"389ecc08",x"70085252",x"70802e8a",x"3884129e",x"cc0c702d",x"ec39810b",x"0b0b0b9e",x"e434833d",x"0d040480",x"3d0d0b0b",x"0b9f9808",x"802e9738",x"0b0b0b0b",x"800b802e",x"8d380b0b",x"0b9f9851",x"0b0b0bf6",x"873f823d",x"0d0404ff",x"3d0d80c4",x"80808452",x"71087082",x"2a708106",x"51515170",x"f338833d",x"0d04ff3d",x"0d80c480",x"80845271",x"0870812a",x"70810651",x"515170f3",x"38738290",x"0a0c833d",x"0d04fe3d",x"0d747080",x"dc808088",x"0c7081ff",x"06ff8311",x"54515371",x"81268d38",x"80fd518a",x"9a2d72a0",x"32518339",x"72518a9a",x"2d843d0d",x"04ff3d0d",x"028f0533",x"5283ffff",x"0b83d00a",x"0c80fe51",x"8a9a2d71",x"518aba2d",x"833d0d04",x"fe3d0d83",x"d00a0870",x"81ff0652",x"528aba2d",x"71882a51",x"8aba2d80",x"fe518a9a",x"2d9efc33",x"81058706",x"52719efc",x"34843d0d",x"04fe3d0d",x"9f803370",x"832b8207",x"81fa0652",x"538ae92d",x"8b882d84",x"3d0d04fe",x"3d0d9f80",x"3370832b",x"810781f9",x"0652538a",x"e92d8b88",x"2d843d0d",x"0482f6ff",x"0b80cc80",x"80880c80",x"0b80cc80",x"80840c9f",x"0b83900a",x"0c04ff3d",x"0d737008",x"515180c8",x"80808470",x"08708480",x"8007720c",x"5252833d",x"0d04ff3d",x"0d80c880",x"80847008",x"70fbffff",x"06720c52",x"52833d0d",x"04a0900b",x"a0800c9e",x"e80ba084",x"0c9b982d",x"ff3d0d73",x"518b710c",x"90115298",x"8080720c",x"80720c70",x"0883ffff",x"06880c83",x"3d0d04fa",x"3d0d787a",x"7dff1e56",x"56585572",x"ff2ea738",x"80568452",x"75750c74",x"0888180c",x"ff125271",x"f3387384",x"15760872",x"0cff1555",x"555272ff",x"2e098106",x"dd38883d",x"0d04f93d",x"0d80d080",x"80845783",x"d00a588c",x"9e2d7651",x"8cc42d9e",x"e8708808",x"84299880",x"84057170",x"8405530c",x"5656fb80",x"84a1ad75",x"0c9ed00b",x"88170c80",x"70780c77",x"0c760870",x"83ffff06",x"515683ff",x"ff780ca0",x"80548808",x"53775276",x"518ce32d",x"76518c82",x"2d770855",x"75752e89",x"3880c351",x"8a9a2dff",x"39a08408",x"5574fba0",x"90ae802e",x"893880c2",x"518a9a2d",x"ff3980d0",x"0a700870",x"ffbf0672",x"0c565689",x"ff2d8cb5",x"2dff3d0d",x"9ef40881",x"119ef40c",x"5183900a",x"700870fe",x"ff06720c",x"5252833d",x"0d04fe3d",x"0d9efc33",x"70832b81",x"80079f80",x"337181f8",x"06075353",x"538ae92d",x"74818007",x"518aba2d",x"8b882d84",x"3d0d04fe",x"3d0d80d0",x"80808453",x"8c9e2d85",x"730c8073",x"0c720870",x"81ff0674",x"5351528c",x"822d7188",x"0c843d0d",x"04fc3d0d",x"76538bb5",x"2d811333",x"82143371",x"81800a29",x"71848080",x"29058316",x"33708280",x"29128418",x"33527105",x"a0800586",x"18851933",x"59525353",x"545654ff",x"135372ff",x"2e913873",x"70810555",x"33527175",x"70810557",x"34e93989",x"518ece2d",x"863d0d04",x"f93d0d79",x"5680d080",x"8084578c",x"9e2d8116",x"33821733",x"71828029",x"05535371",x"802e9438",x"85167255",x"53727081",x"05543377",x"0cff1454",x"73f33883",x"16338417",x"33718280",x"29055652",x"80547375",x"27973873",x"5877770c",x"73167708",x"53537173",x"34811454",x"747426ed",x"3876518c",x"822d9efc",x"3370832b",x"8180079f",x"80337181",x"f8060753",x"53548ae9",x"2d818451",x"8aba2d74",x"882a518a",x"ba2d7451",x"8aba2d80",x"54737527",x"8f387316",x"70335252",x"8aba2d81",x"1454ee39",x"8b882d89",x"3d0d04fc",x"3d0d80d0",x"8080840b",x"81185455",x"8bb52d8c",x"9e2d8675",x"0c74518c",x"822d8c9e",x"2d82750c",x"72708105",x"5433750c",x"72708105",x"5433750c",x"72708105",x"5433750c",x"81ff5472",x"70810554",x"33750cff",x"14547380",x"25f13874",x"518c822d",x"8ef72d88",x"08810652",x"71f63886",x"3d0d04fa",x"3d0d7856",x"80d08080",x"84548c9e",x"2d86740c",x"73518c82",x"2d8c9e2d",x"81ad740c",x"81163382",x"17337182",x"80290583",x"1833760c",x"84183376",x"0c851833",x"760c5852",x"80557477",x"27af3874",x"802e8838",x"8c9e2d81",x"ad740c74",x"16861133",x"750c8711",x"33750c52",x"73518c82",x"2d8ef72d",x"88088106",x"5271f638",x"821555ce",x"398c9e2d",x"84740c73",x"518c822d",x"9efc3370",x"832b8180",x"079f8033",x"7181f806",x"07535353",x"8ae92d81",x"87518aba",x"2d8b882d",x"883d0d04",x"fc3d0d76",x"81113382",x"12337190",x"2b71882b",x"07831433",x"70720788",x"2b841633",x"71075152",x"53565755",x"5288518e",x"ce2d81ff",x"518a9a2d",x"80c48080",x"84547308",x"70812a70",x"81065151",x"5271f338",x"72848080",x"0780c480",x"80840c86",x"3d0d04fd",x"3d0d8ef7",x"2d880888",x"08810653",x"5371f338",x"9efc3370",x"832b8180",x"079f8033",x"7181f806",x"07535354",x"8ae92d81",x"83518aba",x"2d72518a",x"ba2d8b88",x"2d853d0d",x"04fc3d0d",x"800b9ef4",x"0c80709e",x"8c575454",x"74708405",x"56085271",x"802e8a38",x"81138171",x"2b750755",x"52811353",x"8c7327e4",x"38739efc",x"3370832b",x"8180079f",x"80337181",x"f8060754",x"5455538a",x"e92d8181",x"518aba2d",x"9ed05493",x"52737081",x"05553351",x"8aba2dff",x"125271ff",x"2e098106",x"ec387298",x"2a518aba",x"2d72902a",x"518aba2d",x"72882a51",x"8aba2d72",x"518aba2d",x"80518aba",x"2d8f518a",x"ba2d9ec2",x"518aba2d",x"bd84c051",x"8aba2d8b",x"882d863d",x"0d04fe3d",x"0d800b9e",x"f40c9efc",x"3370832b",x"8180079f",x"80337181",x"f8060753",x"53538ae9",x"2d818251",x"8aba2d80",x"d0808084",x"528c9e2d",x"81f90a0b",x"80d08080",x"9c0c7108",x"7252538c",x"822d729f",x"840c7290",x"2a518aba",x"2d9f8408",x"882a518a",x"ba2d9f84",x"08518aba",x"2d8ef72d",x"8808518a",x"ba2d8b88",x"2d843d0d",x"04803d0d",x"810b9ef8",x"0c800b83",x"900a0c85",x"518ece2d",x"823d0d04",x"803d0d80",x"0b9ef80c",x"8be92d86",x"518ece2d",x"823d0d04",x"fd3d0d80",x"d0808084",x"548a518e",x"ce2d8c9e",x"2d9ee874",x"52538cc4",x"2d728808",x"84299880",x"84057170",x"8405530c",x"52fb8084",x"a1ad720c",x"9ed00b88",x"140c7351",x"8c822d89",x"ff2d8cb5",x"2dffb23d",x"0d80d23d",x"0856800b",x"9ef80c80",x"0b9ef40c",x"800bdf80",x"179ed571",x"902a7156",x"56575557",x"72727081",x"05543473",x"882a5372",x"72347382",x"16347598",x"2a52718b",x"16347590",x"2a52718c",x"16347588",x"2a52718d",x"1634758e",x"16348eb1",x"0ba0800c",x"8480b30b",x"80c48080",x"840c80c8",x"8080a453",x"fbffff73",x"08707206",x"750c5354",x"80c88080",x"94700870",x"7606720c",x"5353880b",x"80c08080",x"840c810b",x"900a0c8b",x"e92dfe88",x"880b80dc",x"8080840c",x"81f20b80",x"d00a0c80",x"d0808084",x"7052528c",x"822d8c9e",x"2d71518c",x"822d8c9e",x"2d84720c",x"71518c82",x"2d767756",x"5480c480",x"80840870",x"81065152",x"719e389e",x"f8085372",x"ec389ef4",x"085287e8",x"7227e238",x"72900a0c",x"7283900a",x"0c9b902d",x"82900a08",x"5374802e",x"81d43872",x"80fe2e09",x"8106818d",x"3876802e",x"ffbb3880",x"55827727",x"ffb33883",x"d00a0852",x"71752e09",x"810680c1",x"38883d33",x"70872a81",x"32535371",x"802ea138",x"72870652",x"71ff8e38",x"749f8034",x"749efc34",x"810b9ef8",x"0c748390",x"0a0c8bb5",x"2dfef639",x"72b80670",x"832a9f80",x"33555152",x"71732e87",x"388bcf2d",x"fedf3981",x"13870652",x"719f8034",x"029d0533",x"52718d26",x"fecb3871",x"84299e88",x"0580d13d",x"fde10552",x"70085152",x"712dfeb5",x"397280fd",x"2e098106",x"86388154",x"fea73976",x"829f26a5",x"3873802e",x"87388073",x"a0325454",x"7280dc80",x"80880c80",x"d03d7705",x"fde00552",x"72723481",x"1757fdfd",x"398055fd",x"f8397280",x"fe2e0981",x"06fdee38",x"7457ff0b",x"83d00a0c",x"81775555",x"fddf39ff",x"3d0d9bed",x"2d735280",x"5197992d",x"833d0d04",x"83fffff8",x"0d8d9e04",x"83fffff8",x"0da08804",x"880880c0",x"80808808",x"a080082d",x"50880c81",x"0b900a0c",x"0480700c",x"faad95b4",x"da0b8180",x"8071710c",x"7180082e",x"87387011",x"519bc104",x"519aff2d",x"00000000",x"00000000",x"00000000",x"820b80c0",x"8080900c",x"0b0b0b04",x"0083f00a",x"0b800ba0",x"80721208",x"720c8412",x"5271712e",x"ff05f238",x"028c050d",x"9be00400",x"00000000",x"00000000",x"00000000",x"00fb3d0d",x"77795555",x"80567476",x"25863874",x"30558156",x"73802588",x"38733076",x"81325754",x"80537352",x"745180ca",x"3f880854",x"75802e85",x"38880830",x"5473880c",x"873d0d04",x"fa3d0d78",x"7a575580",x"57747725",x"86387430",x"55815775",x"9f2c5481",x"53757432",x"74315274",x"51943f88",x"08547680",x"2e853888",x"08305473",x"880c883d",x"0d04fc3d",x"0d767853",x"54815380",x"55873971",x"10731054",x"52737226",x"5172802e",x"a7387080",x"2e863871",x"8025e838",x"72802e98",x"38717426",x"89387372",x"31757407",x"56547281",x"2a72812a",x"5353e539",x"73517883",x"38745170",x"880c863d",x"0d04ff3d",x"0d9f8c0b",x"fc055271",x"08ff2e8b",x"38710851",x"702dfc12",x"52f13983",x"3d0d0404",x"ebae3f04",x"00ffffff",x"ff00ffff",x"ffff00ff",x"ffffff00",x"00000a25",x"00000ac2",x"000009eb",x"000007f4",x"00000b2d",x"00000b44",x"000008fb",x"00000998",x"0000079d",x"00000b58",x"0000089b",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000f94",x"02010600",x"00000000",x"05b8d800",x"b4041700",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"ffffffff",x"00000000",x"ffffffff",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000");

begin

  process (clk)
  begin
    if rising_edge(clk) then
      if ENA='1' then
        if WEA='1' then
          RAM(conv_integer(ADDRA) ) := DIA;
        end if;
        DOA <= RAM(conv_integer(ADDRA)) ;
      end if;
    end if;
  end process;  

  process (clk)
  begin
    if rising_edge(clk) then
      if ENB='1' then
        if WEB='1' then
          RAM( conv_integer(ADDRB) ) := DIB;
        end if;
        DOB <= RAM(conv_integer(ADDRB)) ;
      end if;
    end if;
  end process;  
end behave;
