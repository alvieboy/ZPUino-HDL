library IEEE;
use IEEE.std_logic_1164.all; 
use IEEE.std_logic_unsigned.all; 
use ieee.numeric_std.all;

entity bootloader_dp_32 is
  port (
    CLK:              in std_logic;
    WEA:  in std_logic;
    ENA:  in std_logic;
    MASKA:    in std_logic_vector(3 downto 0);
    ADDRA:         in std_logic_vector(11 downto 2);
    DIA:        in std_logic_vector(31 downto 0);
    DOA:         out std_logic_vector(31 downto 0);
    WEB:  in std_logic;
    ENB:  in std_logic;
    ADDRB:         in std_logic_vector(11 downto 2);
    DIB:        in std_logic_vector(31 downto 0);
    MASKB:    in std_logic_vector(3 downto 0);
    DOB:         out std_logic_vector(31 downto 0)
  );
end entity bootloader_dp_32;

architecture behave of bootloader_dp_32 is

  subtype RAM_WORD is STD_LOGIC_VECTOR (31 downto 0);
  type RAM_TABLE is array (0 to 1023) of RAM_WORD;
 shared variable RAM: RAM_TABLE := RAM_TABLE'(
x"0b0b0b97",x"8a040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b97",x"a6040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fd0608",x"72830609",x"81058205",x"832b2a83",x"ffff0652",x"04000000",x"00000000",x"00000000",x"71fd0608",x"83ffff73",x"83060981",x"05820583",x"2b2b0906",x"7383ffff",x"0b0b0b0b",x"83a70400",x"72098105",x"72057373",x"09060906",x"73097306",x"070a8106",x"53510400",x"00000000",x"00000000",x"72722473",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71737109",x"71068106",x"30720a10",x"0a720a10",x"0a31050a",x"81065151",x"53510400",x"00000000",x"72722673",x"732e0753",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"c3040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"720a722b",x"0a535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72729f06",x"0981050b",x"0b0b88a6",x"05040000",x"00000000",x"00000000",x"00000000",x"00000000",x"72722aff",x"739f062a",x"0974090a",x"8106ff05",x"06075351",x"04000000",x"00000000",x"00000000",x"71715351",x"020d0406",x"73830609",x"81058205",x"832b0b2b",x"0772fc06",x"0c515104",x"00000000",x"72098105",x"72050970",x"81050906",x"0a810653",x"51040000",x"00000000",x"00000000",x"00000000",x"72098105",x"72050970",x"81050906",x"0a098106",x"53510400",x"00000000",x"00000000",x"00000000",x"71098105",x"52040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72720981",x"05055351",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097206",x"73730906",x"07535104",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71fc0608",x"72830609",x"81058305",x"1010102a",x"81ff0652",x"04000000",x"00000000",x"00000000",x"71fc0608",x"0b0b0b9c",x"f8738306",x"10100508",x"060b0b0b",x"88a90400",x"00000000",x"00000000",x"0b0b0b88",x"f7040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0b0b0b88",x"df040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"72097081",x"0509060a",x"8106ff05",x"70547106",x"73097274",x"05ff0506",x"07515151",x"04000000",x"72097081",x"0509060a",x"098106ff",x"05705471",x"06730972",x"7405ff05",x"06075151",x"51040000",x"05ff0504",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"810b0b0b",x"0b9dc00c",x"51040000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"71810552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"02840572",x"10100552",x"04000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"717105ff",x"05715351",x"020d0400",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"81d43f94",x"c93f0410",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10101010",x"10105351",x"047381ff",x"06738306",x"09810583",x"05101010",x"2b0772fc",x"060c5151",x"043c0472",x"72807281",x"06ff0509",x"72060571",x"1052720a",x"100a5372",x"ed385151",x"53510488",x"088c0890",x"08757597",x"fc2d5050",x"88085690",x"0c8c0c88",x"0c510488",x"088c0890",x"08757597",x"b82d5050",x"88085690",x"0c8c0c88",x"0c510488",x"088c0890",x"088e812d",x"900c8c0c",x"880c04ff",x"3d0d0b0b",x"0b9dd033",x"5170a638",x"9dcc0870",x"08525270",x"802e9238",x"84129dcc",x"0c702d9d",x"cc087008",x"525270f0",x"38810b0b",x"0b0b9dd0",x"34833d0d",x"0404803d",x"0d0b0b0b",x"9dfc0880",x"2e8e380b",x"0b0b0b80",x"0b802e09",x"81068538",x"823d0d04",x"0b0b0b9d",x"fc510b0b",x"0bf6813f",x"823d0d04",x"04ff3d0d",x"80c48080",x"84527108",x"70822a70",x"81065151",x"5170f338",x"833d0d04",x"ff3d0d80",x"c4808084",x"52710870",x"812a7081",x"06515151",x"70f33873",x"82900a0c",x"833d0d04",x"fe3d0d74",x"7080dc80",x"80880c70",x"81ff06ff",x"83115451",x"53718126",x"8d3880fd",x"518aa02d",x"72a03251",x"83397251",x"8aa02d84",x"3d0d0480",x"3d0d83ff",x"ff0b83d0",x"0a0c80fe",x"518aa02d",x"823d0d04",x"ff3d0d83",x"d00a0870",x"882a5252",x"8ac02d71",x"81ff0651",x"8ac02d80",x"fe518aa0",x"2d833d0d",x"0482f6ff",x"0b80cc80",x"80880c80",x"0b80cc80",x"80840c9f",x"0b83900a",x"0c8e810b",x"a0800c81",x"0b80d00a",x"0c04ff3d",x"0d737008",x"515180c8",x"80808470",x"08708480",x"8007720c",x"5252833d",x"0d04ff3d",x"0d80c880",x"80847008",x"70fbffff",x"06720c52",x"52833d0d",x"04a0900b",x"a0800c9d",x"d40ba084",x"0c979f2d",x"ff3d0d73",x"518b710c",x"90115298",x"8080720c",x"80720c70",x"0883ffff",x"06880c83",x"3d0d04fa",x"3d0d787a",x"7dff1e57",x"57585373",x"ff2ea738",x"80568452",x"75730c72",x"0888180c",x"ff125271",x"f3387484",x"16740872",x"0cff1656",x"565273ff",x"2e098106",x"dd38883d",x"0d04f83d",x"0d80c080",x"80845783",x"d00a598b",x"e62d7651",x"8c8c2d9d",x"d4708808",x"10109880",x"84057170",x"8405530c",x"5656fb80",x"84a1ad75",x"0c9db00b",x"88170c80",x"70780c77",x"0c760883",x"ffff0656",x"9fdf800b",x"88082783",x"38ff3983",x"ffff790c",x"a0805488",x"08537852",x"76518cab",x"2d76518b",x"ca2d7808",x"5574762e",x"893880c3",x"518aa02d",x"ff39a084",x"085574fa",x"a094a680",x"2e893880",x"c2518aa0",x"2dff3990",x"0a700870",x"ffbf0672",x"0c56568a",x"852d8bfd",x"2dff3d0d",x"9de00881",x"119de00c",x"5183900a",x"700870fe",x"ff06720c",x"5252833d",x"0d04803d",x"0d8aef2d",x"72818007",x"518ac02d",x"8b842d82",x"3d0d04fe",x"3d0d80c0",x"80808453",x"8be62d85",x"730c8073",x"0c720870",x"81ff0674",x"5351528b",x"ca2d7188",x"0c843d0d",x"04fc3d0d",x"76811133",x"82123371",x"81800a29",x"71848080",x"29058314",x"33708280",x"29128416",x"33527105",x"a0800586",x"16851733",x"57525353",x"55575553",x"ff135372",x"ff2e9138",x"73708105",x"55335271",x"75708105",x"5734e939",x"89518e9e",x"2d863d0d",x"04f93d0d",x"795780c0",x"80808456",x"8be62d81",x"17338218",x"33718280",x"29055353",x"71802e94",x"38851772",x"55537270",x"81055433",x"760cff14",x"5473f338",x"83173384",x"18337182",x"80290556",x"52805473",x"75279738",x"73587776",x"0c731776",x"08535371",x"73348114",x"54747426",x"ed387551",x"8bca2d8a",x"ef2d8184",x"518ac02d",x"74882a51",x"8ac02d74",x"518ac02d",x"80547375",x"278f3873",x"17703352",x"528ac02d",x"811454ee",x"398b842d",x"893d0d04",x"04fc3d0d",x"76811133",x"82123371",x"902b7188",x"2b078314",x"33707207",x"882b8416",x"33710751",x"52535757",x"54528851",x"8e9e2d81",x"ff518aa0",x"2d80c480",x"80845372",x"0870812a",x"70810651",x"515271f3",x"38738480",x"800780c4",x"8080840c",x"863d0d04",x"fe3d0d8e",x"b32d8808",x"88088106",x"535371f3",x"388aef2d",x"8183518a",x"c02d7251",x"8ac02d8b",x"842d843d",x"0d04fe3d",x"0d800b9d",x"e00c8aef",x"2d818151",x"8ac02d9d",x"b0538f52",x"72708105",x"5433518a",x"c02dff12",x"5271ff2e",x"098106ec",x"388b842d",x"843d0d04",x"fe3d0d80",x"0b9de00c",x"8aef2d81",x"82518ac0",x"2d80c080",x"8084528b",x"e62d81f9",x"0a0b80c0",x"80809c0c",x"71087252",x"538bca2d",x"729de80c",x"72902a51",x"8ac02d9d",x"e808882a",x"518ac02d",x"9de80851",x"8ac02d8e",x"b32d8808",x"518ac02d",x"8b842d84",x"3d0d0480",x"3d0d810b",x"9de40c80",x"0b83900a",x"0c85518e",x"9e2d823d",x"0d04803d",x"0d800b9d",x"e40c8ba5",x"2d86518e",x"9e2d823d",x"0d04fd3d",x"0d80c080",x"8084548a",x"518e9e2d",x"8be62d9d",x"d4745253",x"8c8c2d72",x"88081010",x"98808405",x"71708405",x"530c52fb",x"8084a1ad",x"720c9db0",x"0b88140c",x"73518bca",x"2d8a852d",x"8bfd2dfc",x"3d0d80c0",x"80808470",x"52558bca",x"2d8be62d",x"8b750c76",x"80c08080",x"940c8075",x"0ca08054",x"775383d0",x"0a527451",x"8cab2d74",x"518bca2d",x"8a852d8b",x"fd2dffab",x"3d0d800b",x"9de40c80",x"0b9de00c",x"800b8e81",x"0ba0800c",x"5780c480",x"80845584",x"80b3750c",x"80c88080",x"a453fbff",x"ff730870",x"7206750c",x"535480c8",x"80809470",x"08707606",x"720c5353",x"a87098b4",x"71708405",x"530c9991",x"710c539a",x"aa0b8812",x"0c9bb90b",x"8c120c93",x"af0b9012",x"0c53880b",x"80d08080",x"840c80d0",x"0a538173",x"0c8ba52d",x"8288880b",x"80dc8080",x"840c81f2",x"0b900a0c",x"80c08080",x"84705252",x"8bca2d8b",x"e62d7151",x"8bca2d76",x"77767593",x"3d41415b",x"5b5b83d0",x"0a5c7808",x"70810651",x"52719d38",x"9de40853",x"72f0389d",x"e0085287",x"e87227e6",x"38727e0c",x"7283900a",x"0c97982d",x"82900a08",x"5379802e",x"81b43872",x"80fe2e09",x"810680f4",x"3876802e",x"c138807d",x"7858565a",x"827727ff",x"b53883ff",x"ff7c0c79",x"fe185353",x"79722798",x"3880dc80",x"80887255",x"58721570",x"33790c52",x"81135373",x"7326f238",x"ff167511",x"547505ff",x"05703374",x"33707288",x"2b077f08",x"53515551",x"5271732e",x"098106fe",x"ed387433",x"53728a26",x"fee43872",x"10109d84",x"05755270",x"08515271",x"2dfed339",x"7280fd2e",x"09810686",x"38815bfe",x"c5397682",x"9f269e38",x"7a802e87",x"388073a0",x"32545b80",x"d73d7705",x"fde00552",x"72723481",x"1757fea2",x"39805afe",x"9d397280",x"fe2e0981",x"06fe9338",x"795783ff",x"ff7c0c81",x"775c5afe",x"8539ff3d",x"0d805280",x"5193e62d",x"833d0d04",x"9ffff80d",x"8ce6049f",x"fff80da0",x"88048808",x"8c08a080",x"2d8c0c88",x"0c810b80",x"d00a0c04",x"fb3d0d77",x"79555580",x"56757524",x"ab388074",x"249d3880",x"53735274",x"5180e13f",x"88085475",x"802e8538",x"88083054",x"73880c87",x"3d0d0473",x"30768132",x"5754dc39",x"74305581",x"56738025",x"d238ec39",x"fa3d0d78",x"7a575580",x"57767524",x"a438759f",x"2c548153",x"75743274",x"31527451",x"9b3f8808",x"5476802e",x"85388808",x"30547388",x"0c883d0d",x"04743055",x"8157d739",x"fc3d0d76",x"78535481",x"53807473",x"26525572",x"802e9838",x"70802ea9",x"38807224",x"a4387110",x"73107572",x"26535452",x"72ea3873",x"51788338",x"74517088",x"0c863d0d",x"0472812a",x"72812a53",x"5372802e",x"e6387174",x"26ef3873",x"72317574",x"0774812a",x"74812a55",x"555654e5",x"39fc3d0d",x"7670797b",x"55555555",x"8f72278c",x"38727507",x"83065170",x"802ea738",x"ff125271",x"ff2e9838",x"72708105",x"54337470",x"81055634",x"ff125271",x"ff2e0981",x"06ea3874",x"880c863d",x"0d047451",x"72708405",x"54087170",x"8405530c",x"72708405",x"54087170",x"8405530c",x"72708405",x"54087170",x"8405530c",x"72708405",x"54087170",x"8405530c",x"f0125271",x"8f26c938",x"83722795",x"38727084",x"05540871",x"70840553",x"0cfc1252",x"718326ed",x"387054ff",x"8339fc3d",x"0d767971",x"028c059f",x"05335755",x"53558372",x"278a3874",x"83065170",x"802ea238",x"ff125271",x"ff2e9338",x"73737081",x"055534ff",x"125271ff",x"2e098106",x"ef387488",x"0c863d0d",x"04747488",x"2b750770",x"71902b07",x"5154518f",x"7227a538",x"72717084",x"05530c72",x"71708405",x"530c7271",x"70840553",x"0c727170",x"8405530c",x"f0125271",x"8f26dd38",x"83722790",x"38727170",x"8405530c",x"fc125271",x"8326f238",x"7053ff90",x"39fb3d0d",x"77797072",x"07830653",x"54527093",x"38717373",x"08545654",x"7173082e",x"80c43873",x"75545271",x"337081ff",x"06525470",x"802e9d38",x"72335570",x"752e0981",x"06953881",x"12811471",x"337081ff",x"06545654",x"5270e538",x"72335573",x"81ff0675",x"81ff0671",x"7131880c",x"5252873d",x"0d047109",x"70f7fbfd",x"ff140670",x"f8848281",x"80065151",x"51709738",x"84148416",x"71085456",x"54717508",x"2edc3873",x"755452ff",x"9639800b",x"880c873d",x"0d04ff3d",x"0d9df00b",x"fc057008",x"525270ff",x"2e913870",x"2dfc1270",x"08525270",x"ff2e0981",x"06f13883",x"3d0d0404",x"eca93f04",x"00ffffff",x"ff00ffff",x"ffff00ff",x"ffffff00",x"000008ba",x"000008ec",x"00000894",x"000007ad",x"00000943",x"0000095a",x"00000840",x"00000841",x"00000759",x"0000096e",x"01090600",x"0007ef80",x"05b8d800",x"a4051300",x"00000000",x"00000000",x"00000000",x"00000ef8",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"ffffffff",x"00000000",x"ffffffff",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000");

begin

  process (clk)
  begin
    if rising_edge(clk) then
      if ENA='1' then
        if WEA='1' then
          RAM(conv_integer(ADDRA) ) := DIA;
        end if;
        DOA <= RAM(conv_integer(ADDRA)) ;
      end if;
    end if;
  end process;  

  process (clk)
  begin
    if rising_edge(clk) then
      if ENB='1' then
        if WEB='1' then
          RAM( conv_integer(ADDRB) ) := DIB;
        end if;
        DOB <= RAM(conv_integer(ADDRB)) ;
      end if;
    end if;
  end process;  
end behave;
